-- Tyler Hansen
-- CS232 Final Project
-- genSpriteROM.py
-- generates a ROM file in VHDL from a .ppm image

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity cloud is
port(
X	: in INTEGER RANGE 0 TO 1688;
Y	: in INTEGER RANGE 0 TO 1688;
data : out std_logic_vector (11 downto 0)
);

end entity;

architecture rtl of cloud is
begin
data <=
"000000000000" when X = 0 AND Y = 0 else
"000000000000" when X = 1 AND Y = 0 else
"000000000000" when X = 2 AND Y = 0 else
"000000000000" when X = 3 AND Y = 0 else
"000000000000" when X = 4 AND Y = 0 else
"000000000000" when X = 5 AND Y = 0 else
"000000000000" when X = 6 AND Y = 0 else
"000000000000" when X = 7 AND Y = 0 else
"000000000000" when X = 8 AND Y = 0 else
"000000000000" when X = 9 AND Y = 0 else
"000000000000" when X = 10 AND Y = 0 else
"000000000000" when X = 11 AND Y = 0 else
"000000000000" when X = 12 AND Y = 0 else
"000000000000" when X = 13 AND Y = 0 else
"000000000000" when X = 14 AND Y = 0 else
"000000000000" when X = 15 AND Y = 0 else
"000000000000" when X = 16 AND Y = 0 else
"000000000000" when X = 17 AND Y = 0 else
"000000000000" when X = 18 AND Y = 0 else
"000000000000" when X = 19 AND Y = 0 else
"000000000000" when X = 20 AND Y = 0 else
"000000000000" when X = 21 AND Y = 0 else
"000000000000" when X = 22 AND Y = 0 else
"000000000000" when X = 23 AND Y = 0 else
"000000000000" when X = 24 AND Y = 0 else
"000000000000" when X = 25 AND Y = 0 else
"000000000000" when X = 26 AND Y = 0 else
"000000000000" when X = 27 AND Y = 0 else
"000000000000" when X = 28 AND Y = 0 else
"000000000000" when X = 29 AND Y = 0 else
"000000000000" when X = 30 AND Y = 0 else
"000000000000" when X = 31 AND Y = 0 else
"000000000000" when X = 32 AND Y = 0 else
"000000000000" when X = 33 AND Y = 0 else
"000000000000" when X = 34 AND Y = 0 else
"000000000000" when X = 35 AND Y = 0 else
"000000000000" when X = 36 AND Y = 0 else
"000000000000" when X = 37 AND Y = 0 else
"000000000000" when X = 38 AND Y = 0 else
"000000000000" when X = 39 AND Y = 0 else
"000000000000" when X = 40 AND Y = 0 else
"000000000000" when X = 41 AND Y = 0 else
"000000000000" when X = 42 AND Y = 0 else
"000000000000" when X = 43 AND Y = 0 else
"000000000000" when X = 44 AND Y = 0 else
"000000000000" when X = 45 AND Y = 0 else
"000000000000" when X = 46 AND Y = 0 else
"000000000000" when X = 47 AND Y = 0 else
"000000000000" when X = 48 AND Y = 0 else
"000000000000" when X = 49 AND Y = 0 else
"000000000000" when X = 50 AND Y = 0 else
"000000000000" when X = 51 AND Y = 0 else
"000000000000" when X = 52 AND Y = 0 else
"000000000000" when X = 53 AND Y = 0 else
"000000000000" when X = 54 AND Y = 0 else
"000000000000" when X = 55 AND Y = 0 else
"000000000000" when X = 56 AND Y = 0 else
"000000000000" when X = 57 AND Y = 0 else
"000000000000" when X = 58 AND Y = 0 else
"000000000000" when X = 59 AND Y = 0 else
"000000000000" when X = 60 AND Y = 0 else
"000000000000" when X = 61 AND Y = 0 else
"000000000000" when X = 62 AND Y = 0 else
"000000000000" when X = 63 AND Y = 0 else
"000000000000" when X = 64 AND Y = 0 else
"000000000000" when X = 65 AND Y = 0 else
"000000000000" when X = 66 AND Y = 0 else
"000000000000" when X = 67 AND Y = 0 else
"000000000000" when X = 68 AND Y = 0 else
"000000000000" when X = 69 AND Y = 0 else
"000000000000" when X = 70 AND Y = 0 else
"000000000000" when X = 71 AND Y = 0 else
"000000000000" when X = 72 AND Y = 0 else
"000000000000" when X = 73 AND Y = 0 else
"000000000000" when X = 74 AND Y = 0 else
"000000000000" when X = 75 AND Y = 0 else
"000000000000" when X = 76 AND Y = 0 else
"000000000000" when X = 77 AND Y = 0 else
"000000000000" when X = 78 AND Y = 0 else
"000000000000" when X = 79 AND Y = 0 else
"111111111111" when X = 80 AND Y = 0 else
"111111111111" when X = 81 AND Y = 0 else
"111111111111" when X = 82 AND Y = 0 else
"111111111111" when X = 83 AND Y = 0 else
"111111111111" when X = 84 AND Y = 0 else
"111111111111" when X = 85 AND Y = 0 else
"111111111111" when X = 86 AND Y = 0 else
"111111111111" when X = 87 AND Y = 0 else
"111111111111" when X = 88 AND Y = 0 else
"111111111111" when X = 89 AND Y = 0 else
"111111111111" when X = 90 AND Y = 0 else
"111111111111" when X = 91 AND Y = 0 else
"111111111111" when X = 92 AND Y = 0 else
"111111111111" when X = 93 AND Y = 0 else
"111111111111" when X = 94 AND Y = 0 else
"111111111111" when X = 95 AND Y = 0 else
"111111111111" when X = 96 AND Y = 0 else
"111111111111" when X = 97 AND Y = 0 else
"111111111111" when X = 98 AND Y = 0 else
"111111111111" when X = 99 AND Y = 0 else
"111111111111" when X = 100 AND Y = 0 else
"111111111111" when X = 101 AND Y = 0 else
"111111111111" when X = 102 AND Y = 0 else
"111111111111" when X = 103 AND Y = 0 else
"111111111111" when X = 104 AND Y = 0 else
"111111111111" when X = 105 AND Y = 0 else
"111111111111" when X = 106 AND Y = 0 else
"111111111111" when X = 107 AND Y = 0 else
"111111111111" when X = 108 AND Y = 0 else
"111111111111" when X = 109 AND Y = 0 else
"111111111111" when X = 110 AND Y = 0 else
"111111111111" when X = 111 AND Y = 0 else
"111111111111" when X = 112 AND Y = 0 else
"111111111111" when X = 113 AND Y = 0 else
"111111111111" when X = 114 AND Y = 0 else
"111111111111" when X = 115 AND Y = 0 else
"111111111111" when X = 116 AND Y = 0 else
"111111111111" when X = 117 AND Y = 0 else
"111111111111" when X = 118 AND Y = 0 else
"111111111111" when X = 119 AND Y = 0 else
"111111111111" when X = 120 AND Y = 0 else
"111111111111" when X = 121 AND Y = 0 else
"111111111111" when X = 122 AND Y = 0 else
"111111111111" when X = 123 AND Y = 0 else
"111111111111" when X = 124 AND Y = 0 else
"111111111111" when X = 125 AND Y = 0 else
"111111111111" when X = 126 AND Y = 0 else
"111111111111" when X = 127 AND Y = 0 else
"111111111111" when X = 128 AND Y = 0 else
"111111111111" when X = 129 AND Y = 0 else
"111111111111" when X = 130 AND Y = 0 else
"111111111111" when X = 131 AND Y = 0 else
"111111111111" when X = 132 AND Y = 0 else
"111111111111" when X = 133 AND Y = 0 else
"111111111111" when X = 134 AND Y = 0 else
"111111111111" when X = 135 AND Y = 0 else
"111111111111" when X = 136 AND Y = 0 else
"111111111111" when X = 137 AND Y = 0 else
"111111111111" when X = 138 AND Y = 0 else
"111111111111" when X = 139 AND Y = 0 else
"000000000000" when X = 140 AND Y = 0 else
"000000000000" when X = 141 AND Y = 0 else
"000000000000" when X = 142 AND Y = 0 else
"000000000000" when X = 143 AND Y = 0 else
"000000000000" when X = 144 AND Y = 0 else
"000000000000" when X = 145 AND Y = 0 else
"000000000000" when X = 146 AND Y = 0 else
"000000000000" when X = 147 AND Y = 0 else
"000000000000" when X = 148 AND Y = 0 else
"000000000000" when X = 149 AND Y = 0 else
"000000000000" when X = 150 AND Y = 0 else
"000000000000" when X = 151 AND Y = 0 else
"000000000000" when X = 152 AND Y = 0 else
"000000000000" when X = 153 AND Y = 0 else
"000000000000" when X = 154 AND Y = 0 else
"000000000000" when X = 155 AND Y = 0 else
"000000000000" when X = 156 AND Y = 0 else
"000000000000" when X = 157 AND Y = 0 else
"000000000000" when X = 158 AND Y = 0 else
"000000000000" when X = 159 AND Y = 0 else
"000000000000" when X = 160 AND Y = 0 else
"000000000000" when X = 161 AND Y = 0 else
"000000000000" when X = 162 AND Y = 0 else
"000000000000" when X = 163 AND Y = 0 else
"000000000000" when X = 164 AND Y = 0 else
"000000000000" when X = 165 AND Y = 0 else
"000000000000" when X = 166 AND Y = 0 else
"000000000000" when X = 167 AND Y = 0 else
"000000000000" when X = 168 AND Y = 0 else
"000000000000" when X = 169 AND Y = 0 else
"000000000000" when X = 170 AND Y = 0 else
"000000000000" when X = 171 AND Y = 0 else
"000000000000" when X = 172 AND Y = 0 else
"000000000000" when X = 173 AND Y = 0 else
"000000000000" when X = 174 AND Y = 0 else
"000000000000" when X = 175 AND Y = 0 else
"000000000000" when X = 176 AND Y = 0 else
"000000000000" when X = 177 AND Y = 0 else
"000000000000" when X = 178 AND Y = 0 else
"000000000000" when X = 179 AND Y = 0 else
"000000000000" when X = 180 AND Y = 0 else
"000000000000" when X = 181 AND Y = 0 else
"000000000000" when X = 182 AND Y = 0 else
"000000000000" when X = 183 AND Y = 0 else
"000000000000" when X = 184 AND Y = 0 else
"000000000000" when X = 185 AND Y = 0 else
"000000000000" when X = 186 AND Y = 0 else
"000000000000" when X = 187 AND Y = 0 else
"000000000000" when X = 188 AND Y = 0 else
"000000000000" when X = 189 AND Y = 0 else
"000000000000" when X = 190 AND Y = 0 else
"000000000000" when X = 191 AND Y = 0 else
"000000000000" when X = 192 AND Y = 0 else
"000000000000" when X = 193 AND Y = 0 else
"000000000000" when X = 194 AND Y = 0 else
"000000000000" when X = 195 AND Y = 0 else
"000000000000" when X = 196 AND Y = 0 else
"000000000000" when X = 197 AND Y = 0 else
"000000000000" when X = 198 AND Y = 0 else
"000000000000" when X = 199 AND Y = 0 else
"000000000000" when X = 200 AND Y = 0 else
"000000000000" when X = 201 AND Y = 0 else
"000000000000" when X = 202 AND Y = 0 else
"000000000000" when X = 203 AND Y = 0 else
"000000000000" when X = 204 AND Y = 0 else
"000000000000" when X = 205 AND Y = 0 else
"000000000000" when X = 206 AND Y = 0 else
"000000000000" when X = 207 AND Y = 0 else
"000000000000" when X = 208 AND Y = 0 else
"000000000000" when X = 209 AND Y = 0 else
"000000000000" when X = 210 AND Y = 0 else
"000000000000" when X = 211 AND Y = 0 else
"000000000000" when X = 212 AND Y = 0 else
"000000000000" when X = 213 AND Y = 0 else
"000000000000" when X = 214 AND Y = 0 else
"000000000000" when X = 215 AND Y = 0 else
"000000000000" when X = 216 AND Y = 0 else
"000000000000" when X = 217 AND Y = 0 else
"000000000000" when X = 218 AND Y = 0 else
"000000000000" when X = 219 AND Y = 0 else
"000000000000" when X = 220 AND Y = 0 else
"000000000000" when X = 221 AND Y = 0 else
"000000000000" when X = 222 AND Y = 0 else
"000000000000" when X = 223 AND Y = 0 else
"000000000000" when X = 224 AND Y = 0 else
"000000000000" when X = 225 AND Y = 0 else
"000000000000" when X = 226 AND Y = 0 else
"000000000000" when X = 227 AND Y = 0 else
"000000000000" when X = 228 AND Y = 0 else
"000000000000" when X = 229 AND Y = 0 else
"000000000000" when X = 230 AND Y = 0 else
"000000000000" when X = 231 AND Y = 0 else
"000000000000" when X = 232 AND Y = 0 else
"000000000000" when X = 233 AND Y = 0 else
"000000000000" when X = 234 AND Y = 0 else
"000000000000" when X = 235 AND Y = 0 else
"000000000000" when X = 236 AND Y = 0 else
"000000000000" when X = 237 AND Y = 0 else
"000000000000" when X = 238 AND Y = 0 else
"000000000000" when X = 239 AND Y = 0 else
"000000000000" when X = 240 AND Y = 0 else
"000000000000" when X = 241 AND Y = 0 else
"000000000000" when X = 242 AND Y = 0 else
"000000000000" when X = 243 AND Y = 0 else
"000000000000" when X = 244 AND Y = 0 else
"000000000000" when X = 245 AND Y = 0 else
"000000000000" when X = 246 AND Y = 0 else
"000000000000" when X = 247 AND Y = 0 else
"000000000000" when X = 248 AND Y = 0 else
"000000000000" when X = 249 AND Y = 0 else
"000000000000" when X = 250 AND Y = 0 else
"000000000000" when X = 251 AND Y = 0 else
"000000000000" when X = 252 AND Y = 0 else
"000000000000" when X = 253 AND Y = 0 else
"000000000000" when X = 254 AND Y = 0 else
"000000000000" when X = 255 AND Y = 0 else
"000000000000" when X = 256 AND Y = 0 else
"000000000000" when X = 257 AND Y = 0 else
"000000000000" when X = 258 AND Y = 0 else
"000000000000" when X = 259 AND Y = 0 else
"000000000000" when X = 260 AND Y = 0 else
"000000000000" when X = 261 AND Y = 0 else
"000000000000" when X = 262 AND Y = 0 else
"000000000000" when X = 263 AND Y = 0 else
"000000000000" when X = 264 AND Y = 0 else
"000000000000" when X = 265 AND Y = 0 else
"000000000000" when X = 266 AND Y = 0 else
"000000000000" when X = 267 AND Y = 0 else
"000000000000" when X = 268 AND Y = 0 else
"000000000000" when X = 269 AND Y = 0 else
"000000000000" when X = 270 AND Y = 0 else
"000000000000" when X = 271 AND Y = 0 else
"000000000000" when X = 272 AND Y = 0 else
"000000000000" when X = 273 AND Y = 0 else
"000000000000" when X = 274 AND Y = 0 else
"000000000000" when X = 275 AND Y = 0 else
"000000000000" when X = 276 AND Y = 0 else
"000000000000" when X = 277 AND Y = 0 else
"000000000000" when X = 278 AND Y = 0 else
"000000000000" when X = 279 AND Y = 0 else
"000000000000" when X = 280 AND Y = 0 else
"000000000000" when X = 281 AND Y = 0 else
"000000000000" when X = 282 AND Y = 0 else
"000000000000" when X = 283 AND Y = 0 else
"000000000000" when X = 284 AND Y = 0 else
"000000000000" when X = 285 AND Y = 0 else
"000000000000" when X = 286 AND Y = 0 else
"000000000000" when X = 287 AND Y = 0 else
"000000000000" when X = 288 AND Y = 0 else
"000000000000" when X = 289 AND Y = 0 else
"000000000000" when X = 290 AND Y = 0 else
"000000000000" when X = 291 AND Y = 0 else
"000000000000" when X = 292 AND Y = 0 else
"000000000000" when X = 293 AND Y = 0 else
"000000000000" when X = 294 AND Y = 0 else
"000000000000" when X = 295 AND Y = 0 else
"000000000000" when X = 296 AND Y = 0 else
"000000000000" when X = 297 AND Y = 0 else
"000000000000" when X = 298 AND Y = 0 else
"000000000000" when X = 299 AND Y = 0 else
"000000000000" when X = 300 AND Y = 0 else
"000000000000" when X = 301 AND Y = 0 else
"000000000000" when X = 302 AND Y = 0 else
"000000000000" when X = 303 AND Y = 0 else
"000000000000" when X = 304 AND Y = 0 else
"000000000000" when X = 305 AND Y = 0 else
"000000000000" when X = 306 AND Y = 0 else
"000000000000" when X = 307 AND Y = 0 else
"000000000000" when X = 308 AND Y = 0 else
"000000000000" when X = 309 AND Y = 0 else
"000000000000" when X = 310 AND Y = 0 else
"000000000000" when X = 311 AND Y = 0 else
"000000000000" when X = 312 AND Y = 0 else
"000000000000" when X = 313 AND Y = 0 else
"000000000000" when X = 314 AND Y = 0 else
"000000000000" when X = 315 AND Y = 0 else
"000000000000" when X = 316 AND Y = 0 else
"000000000000" when X = 317 AND Y = 0 else
"000000000000" when X = 318 AND Y = 0 else
"000000000000" when X = 319 AND Y = 0 else
"000000000000" when X = 320 AND Y = 0 else
"000000000000" when X = 321 AND Y = 0 else
"000000000000" when X = 322 AND Y = 0 else
"000000000000" when X = 323 AND Y = 0 else
"000000000000" when X = 324 AND Y = 0 else
"000000000000" when X = 0 AND Y = 1 else
"000000000000" when X = 1 AND Y = 1 else
"000000000000" when X = 2 AND Y = 1 else
"000000000000" when X = 3 AND Y = 1 else
"000000000000" when X = 4 AND Y = 1 else
"000000000000" when X = 5 AND Y = 1 else
"000000000000" when X = 6 AND Y = 1 else
"000000000000" when X = 7 AND Y = 1 else
"000000000000" when X = 8 AND Y = 1 else
"000000000000" when X = 9 AND Y = 1 else
"000000000000" when X = 10 AND Y = 1 else
"000000000000" when X = 11 AND Y = 1 else
"000000000000" when X = 12 AND Y = 1 else
"000000000000" when X = 13 AND Y = 1 else
"000000000000" when X = 14 AND Y = 1 else
"000000000000" when X = 15 AND Y = 1 else
"000000000000" when X = 16 AND Y = 1 else
"000000000000" when X = 17 AND Y = 1 else
"000000000000" when X = 18 AND Y = 1 else
"000000000000" when X = 19 AND Y = 1 else
"000000000000" when X = 20 AND Y = 1 else
"000000000000" when X = 21 AND Y = 1 else
"000000000000" when X = 22 AND Y = 1 else
"000000000000" when X = 23 AND Y = 1 else
"000000000000" when X = 24 AND Y = 1 else
"000000000000" when X = 25 AND Y = 1 else
"000000000000" when X = 26 AND Y = 1 else
"000000000000" when X = 27 AND Y = 1 else
"000000000000" when X = 28 AND Y = 1 else
"000000000000" when X = 29 AND Y = 1 else
"000000000000" when X = 30 AND Y = 1 else
"000000000000" when X = 31 AND Y = 1 else
"000000000000" when X = 32 AND Y = 1 else
"000000000000" when X = 33 AND Y = 1 else
"000000000000" when X = 34 AND Y = 1 else
"000000000000" when X = 35 AND Y = 1 else
"000000000000" when X = 36 AND Y = 1 else
"000000000000" when X = 37 AND Y = 1 else
"000000000000" when X = 38 AND Y = 1 else
"000000000000" when X = 39 AND Y = 1 else
"000000000000" when X = 40 AND Y = 1 else
"000000000000" when X = 41 AND Y = 1 else
"000000000000" when X = 42 AND Y = 1 else
"000000000000" when X = 43 AND Y = 1 else
"000000000000" when X = 44 AND Y = 1 else
"000000000000" when X = 45 AND Y = 1 else
"000000000000" when X = 46 AND Y = 1 else
"000000000000" when X = 47 AND Y = 1 else
"000000000000" when X = 48 AND Y = 1 else
"000000000000" when X = 49 AND Y = 1 else
"000000000000" when X = 50 AND Y = 1 else
"000000000000" when X = 51 AND Y = 1 else
"000000000000" when X = 52 AND Y = 1 else
"000000000000" when X = 53 AND Y = 1 else
"000000000000" when X = 54 AND Y = 1 else
"000000000000" when X = 55 AND Y = 1 else
"000000000000" when X = 56 AND Y = 1 else
"000000000000" when X = 57 AND Y = 1 else
"000000000000" when X = 58 AND Y = 1 else
"000000000000" when X = 59 AND Y = 1 else
"000000000000" when X = 60 AND Y = 1 else
"000000000000" when X = 61 AND Y = 1 else
"000000000000" when X = 62 AND Y = 1 else
"000000000000" when X = 63 AND Y = 1 else
"000000000000" when X = 64 AND Y = 1 else
"000000000000" when X = 65 AND Y = 1 else
"000000000000" when X = 66 AND Y = 1 else
"000000000000" when X = 67 AND Y = 1 else
"000000000000" when X = 68 AND Y = 1 else
"000000000000" when X = 69 AND Y = 1 else
"000000000000" when X = 70 AND Y = 1 else
"000000000000" when X = 71 AND Y = 1 else
"000000000000" when X = 72 AND Y = 1 else
"000000000000" when X = 73 AND Y = 1 else
"000000000000" when X = 74 AND Y = 1 else
"000000000000" when X = 75 AND Y = 1 else
"000000000000" when X = 76 AND Y = 1 else
"000000000000" when X = 77 AND Y = 1 else
"000000000000" when X = 78 AND Y = 1 else
"000000000000" when X = 79 AND Y = 1 else
"111111111111" when X = 80 AND Y = 1 else
"111111111111" when X = 81 AND Y = 1 else
"111111111111" when X = 82 AND Y = 1 else
"111111111111" when X = 83 AND Y = 1 else
"111111111111" when X = 84 AND Y = 1 else
"111111111111" when X = 85 AND Y = 1 else
"111111111111" when X = 86 AND Y = 1 else
"111111111111" when X = 87 AND Y = 1 else
"111111111111" when X = 88 AND Y = 1 else
"111111111111" when X = 89 AND Y = 1 else
"111111111111" when X = 90 AND Y = 1 else
"111111111111" when X = 91 AND Y = 1 else
"111111111111" when X = 92 AND Y = 1 else
"111111111111" when X = 93 AND Y = 1 else
"111111111111" when X = 94 AND Y = 1 else
"111111111111" when X = 95 AND Y = 1 else
"111111111111" when X = 96 AND Y = 1 else
"111111111111" when X = 97 AND Y = 1 else
"111111111111" when X = 98 AND Y = 1 else
"111111111111" when X = 99 AND Y = 1 else
"111111111111" when X = 100 AND Y = 1 else
"111111111111" when X = 101 AND Y = 1 else
"111111111111" when X = 102 AND Y = 1 else
"111111111111" when X = 103 AND Y = 1 else
"111111111111" when X = 104 AND Y = 1 else
"111111111111" when X = 105 AND Y = 1 else
"111111111111" when X = 106 AND Y = 1 else
"111111111111" when X = 107 AND Y = 1 else
"111111111111" when X = 108 AND Y = 1 else
"111111111111" when X = 109 AND Y = 1 else
"111111111111" when X = 110 AND Y = 1 else
"111111111111" when X = 111 AND Y = 1 else
"111111111111" when X = 112 AND Y = 1 else
"111111111111" when X = 113 AND Y = 1 else
"111111111111" when X = 114 AND Y = 1 else
"111111111111" when X = 115 AND Y = 1 else
"111111111111" when X = 116 AND Y = 1 else
"111111111111" when X = 117 AND Y = 1 else
"111111111111" when X = 118 AND Y = 1 else
"111111111111" when X = 119 AND Y = 1 else
"111111111111" when X = 120 AND Y = 1 else
"111111111111" when X = 121 AND Y = 1 else
"111111111111" when X = 122 AND Y = 1 else
"111111111111" when X = 123 AND Y = 1 else
"111111111111" when X = 124 AND Y = 1 else
"111111111111" when X = 125 AND Y = 1 else
"111111111111" when X = 126 AND Y = 1 else
"111111111111" when X = 127 AND Y = 1 else
"111111111111" when X = 128 AND Y = 1 else
"111111111111" when X = 129 AND Y = 1 else
"111111111111" when X = 130 AND Y = 1 else
"111111111111" when X = 131 AND Y = 1 else
"111111111111" when X = 132 AND Y = 1 else
"111111111111" when X = 133 AND Y = 1 else
"111111111111" when X = 134 AND Y = 1 else
"111111111111" when X = 135 AND Y = 1 else
"111111111111" when X = 136 AND Y = 1 else
"111111111111" when X = 137 AND Y = 1 else
"111111111111" when X = 138 AND Y = 1 else
"111111111111" when X = 139 AND Y = 1 else
"000000000000" when X = 140 AND Y = 1 else
"000000000000" when X = 141 AND Y = 1 else
"000000000000" when X = 142 AND Y = 1 else
"000000000000" when X = 143 AND Y = 1 else
"000000000000" when X = 144 AND Y = 1 else
"000000000000" when X = 145 AND Y = 1 else
"000000000000" when X = 146 AND Y = 1 else
"000000000000" when X = 147 AND Y = 1 else
"000000000000" when X = 148 AND Y = 1 else
"000000000000" when X = 149 AND Y = 1 else
"000000000000" when X = 150 AND Y = 1 else
"000000000000" when X = 151 AND Y = 1 else
"000000000000" when X = 152 AND Y = 1 else
"000000000000" when X = 153 AND Y = 1 else
"000000000000" when X = 154 AND Y = 1 else
"000000000000" when X = 155 AND Y = 1 else
"000000000000" when X = 156 AND Y = 1 else
"000000000000" when X = 157 AND Y = 1 else
"000000000000" when X = 158 AND Y = 1 else
"000000000000" when X = 159 AND Y = 1 else
"000000000000" when X = 160 AND Y = 1 else
"000000000000" when X = 161 AND Y = 1 else
"000000000000" when X = 162 AND Y = 1 else
"000000000000" when X = 163 AND Y = 1 else
"000000000000" when X = 164 AND Y = 1 else
"000000000000" when X = 165 AND Y = 1 else
"000000000000" when X = 166 AND Y = 1 else
"000000000000" when X = 167 AND Y = 1 else
"000000000000" when X = 168 AND Y = 1 else
"000000000000" when X = 169 AND Y = 1 else
"000000000000" when X = 170 AND Y = 1 else
"000000000000" when X = 171 AND Y = 1 else
"000000000000" when X = 172 AND Y = 1 else
"000000000000" when X = 173 AND Y = 1 else
"000000000000" when X = 174 AND Y = 1 else
"000000000000" when X = 175 AND Y = 1 else
"000000000000" when X = 176 AND Y = 1 else
"000000000000" when X = 177 AND Y = 1 else
"000000000000" when X = 178 AND Y = 1 else
"000000000000" when X = 179 AND Y = 1 else
"000000000000" when X = 180 AND Y = 1 else
"000000000000" when X = 181 AND Y = 1 else
"000000000000" when X = 182 AND Y = 1 else
"000000000000" when X = 183 AND Y = 1 else
"000000000000" when X = 184 AND Y = 1 else
"000000000000" when X = 185 AND Y = 1 else
"000000000000" when X = 186 AND Y = 1 else
"000000000000" when X = 187 AND Y = 1 else
"000000000000" when X = 188 AND Y = 1 else
"000000000000" when X = 189 AND Y = 1 else
"000000000000" when X = 190 AND Y = 1 else
"000000000000" when X = 191 AND Y = 1 else
"000000000000" when X = 192 AND Y = 1 else
"000000000000" when X = 193 AND Y = 1 else
"000000000000" when X = 194 AND Y = 1 else
"000000000000" when X = 195 AND Y = 1 else
"000000000000" when X = 196 AND Y = 1 else
"000000000000" when X = 197 AND Y = 1 else
"000000000000" when X = 198 AND Y = 1 else
"000000000000" when X = 199 AND Y = 1 else
"000000000000" when X = 200 AND Y = 1 else
"000000000000" when X = 201 AND Y = 1 else
"000000000000" when X = 202 AND Y = 1 else
"000000000000" when X = 203 AND Y = 1 else
"000000000000" when X = 204 AND Y = 1 else
"000000000000" when X = 205 AND Y = 1 else
"000000000000" when X = 206 AND Y = 1 else
"000000000000" when X = 207 AND Y = 1 else
"000000000000" when X = 208 AND Y = 1 else
"000000000000" when X = 209 AND Y = 1 else
"000000000000" when X = 210 AND Y = 1 else
"000000000000" when X = 211 AND Y = 1 else
"000000000000" when X = 212 AND Y = 1 else
"000000000000" when X = 213 AND Y = 1 else
"000000000000" when X = 214 AND Y = 1 else
"000000000000" when X = 215 AND Y = 1 else
"000000000000" when X = 216 AND Y = 1 else
"000000000000" when X = 217 AND Y = 1 else
"000000000000" when X = 218 AND Y = 1 else
"000000000000" when X = 219 AND Y = 1 else
"000000000000" when X = 220 AND Y = 1 else
"000000000000" when X = 221 AND Y = 1 else
"000000000000" when X = 222 AND Y = 1 else
"000000000000" when X = 223 AND Y = 1 else
"000000000000" when X = 224 AND Y = 1 else
"000000000000" when X = 225 AND Y = 1 else
"000000000000" when X = 226 AND Y = 1 else
"000000000000" when X = 227 AND Y = 1 else
"000000000000" when X = 228 AND Y = 1 else
"000000000000" when X = 229 AND Y = 1 else
"000000000000" when X = 230 AND Y = 1 else
"000000000000" when X = 231 AND Y = 1 else
"000000000000" when X = 232 AND Y = 1 else
"000000000000" when X = 233 AND Y = 1 else
"000000000000" when X = 234 AND Y = 1 else
"000000000000" when X = 235 AND Y = 1 else
"000000000000" when X = 236 AND Y = 1 else
"000000000000" when X = 237 AND Y = 1 else
"000000000000" when X = 238 AND Y = 1 else
"000000000000" when X = 239 AND Y = 1 else
"000000000000" when X = 240 AND Y = 1 else
"000000000000" when X = 241 AND Y = 1 else
"000000000000" when X = 242 AND Y = 1 else
"000000000000" when X = 243 AND Y = 1 else
"000000000000" when X = 244 AND Y = 1 else
"000000000000" when X = 245 AND Y = 1 else
"000000000000" when X = 246 AND Y = 1 else
"000000000000" when X = 247 AND Y = 1 else
"000000000000" when X = 248 AND Y = 1 else
"000000000000" when X = 249 AND Y = 1 else
"000000000000" when X = 250 AND Y = 1 else
"000000000000" when X = 251 AND Y = 1 else
"000000000000" when X = 252 AND Y = 1 else
"000000000000" when X = 253 AND Y = 1 else
"000000000000" when X = 254 AND Y = 1 else
"000000000000" when X = 255 AND Y = 1 else
"000000000000" when X = 256 AND Y = 1 else
"000000000000" when X = 257 AND Y = 1 else
"000000000000" when X = 258 AND Y = 1 else
"000000000000" when X = 259 AND Y = 1 else
"000000000000" when X = 260 AND Y = 1 else
"000000000000" when X = 261 AND Y = 1 else
"000000000000" when X = 262 AND Y = 1 else
"000000000000" when X = 263 AND Y = 1 else
"000000000000" when X = 264 AND Y = 1 else
"000000000000" when X = 265 AND Y = 1 else
"000000000000" when X = 266 AND Y = 1 else
"000000000000" when X = 267 AND Y = 1 else
"000000000000" when X = 268 AND Y = 1 else
"000000000000" when X = 269 AND Y = 1 else
"000000000000" when X = 270 AND Y = 1 else
"000000000000" when X = 271 AND Y = 1 else
"000000000000" when X = 272 AND Y = 1 else
"000000000000" when X = 273 AND Y = 1 else
"000000000000" when X = 274 AND Y = 1 else
"000000000000" when X = 275 AND Y = 1 else
"000000000000" when X = 276 AND Y = 1 else
"000000000000" when X = 277 AND Y = 1 else
"000000000000" when X = 278 AND Y = 1 else
"000000000000" when X = 279 AND Y = 1 else
"000000000000" when X = 280 AND Y = 1 else
"000000000000" when X = 281 AND Y = 1 else
"000000000000" when X = 282 AND Y = 1 else
"000000000000" when X = 283 AND Y = 1 else
"000000000000" when X = 284 AND Y = 1 else
"000000000000" when X = 285 AND Y = 1 else
"000000000000" when X = 286 AND Y = 1 else
"000000000000" when X = 287 AND Y = 1 else
"000000000000" when X = 288 AND Y = 1 else
"000000000000" when X = 289 AND Y = 1 else
"000000000000" when X = 290 AND Y = 1 else
"000000000000" when X = 291 AND Y = 1 else
"000000000000" when X = 292 AND Y = 1 else
"000000000000" when X = 293 AND Y = 1 else
"000000000000" when X = 294 AND Y = 1 else
"000000000000" when X = 295 AND Y = 1 else
"000000000000" when X = 296 AND Y = 1 else
"000000000000" when X = 297 AND Y = 1 else
"000000000000" when X = 298 AND Y = 1 else
"000000000000" when X = 299 AND Y = 1 else
"000000000000" when X = 300 AND Y = 1 else
"000000000000" when X = 301 AND Y = 1 else
"000000000000" when X = 302 AND Y = 1 else
"000000000000" when X = 303 AND Y = 1 else
"000000000000" when X = 304 AND Y = 1 else
"000000000000" when X = 305 AND Y = 1 else
"000000000000" when X = 306 AND Y = 1 else
"000000000000" when X = 307 AND Y = 1 else
"000000000000" when X = 308 AND Y = 1 else
"000000000000" when X = 309 AND Y = 1 else
"000000000000" when X = 310 AND Y = 1 else
"000000000000" when X = 311 AND Y = 1 else
"000000000000" when X = 312 AND Y = 1 else
"000000000000" when X = 313 AND Y = 1 else
"000000000000" when X = 314 AND Y = 1 else
"000000000000" when X = 315 AND Y = 1 else
"000000000000" when X = 316 AND Y = 1 else
"000000000000" when X = 317 AND Y = 1 else
"000000000000" when X = 318 AND Y = 1 else
"000000000000" when X = 319 AND Y = 1 else
"000000000000" when X = 320 AND Y = 1 else
"000000000000" when X = 321 AND Y = 1 else
"000000000000" when X = 322 AND Y = 1 else
"000000000000" when X = 323 AND Y = 1 else
"000000000000" when X = 324 AND Y = 1 else
"000000000000" when X = 0 AND Y = 2 else
"000000000000" when X = 1 AND Y = 2 else
"000000000000" when X = 2 AND Y = 2 else
"000000000000" when X = 3 AND Y = 2 else
"000000000000" when X = 4 AND Y = 2 else
"000000000000" when X = 5 AND Y = 2 else
"000000000000" when X = 6 AND Y = 2 else
"000000000000" when X = 7 AND Y = 2 else
"000000000000" when X = 8 AND Y = 2 else
"000000000000" when X = 9 AND Y = 2 else
"000000000000" when X = 10 AND Y = 2 else
"000000000000" when X = 11 AND Y = 2 else
"000000000000" when X = 12 AND Y = 2 else
"000000000000" when X = 13 AND Y = 2 else
"000000000000" when X = 14 AND Y = 2 else
"000000000000" when X = 15 AND Y = 2 else
"000000000000" when X = 16 AND Y = 2 else
"000000000000" when X = 17 AND Y = 2 else
"000000000000" when X = 18 AND Y = 2 else
"000000000000" when X = 19 AND Y = 2 else
"000000000000" when X = 20 AND Y = 2 else
"000000000000" when X = 21 AND Y = 2 else
"000000000000" when X = 22 AND Y = 2 else
"000000000000" when X = 23 AND Y = 2 else
"000000000000" when X = 24 AND Y = 2 else
"000000000000" when X = 25 AND Y = 2 else
"000000000000" when X = 26 AND Y = 2 else
"000000000000" when X = 27 AND Y = 2 else
"000000000000" when X = 28 AND Y = 2 else
"000000000000" when X = 29 AND Y = 2 else
"000000000000" when X = 30 AND Y = 2 else
"000000000000" when X = 31 AND Y = 2 else
"000000000000" when X = 32 AND Y = 2 else
"000000000000" when X = 33 AND Y = 2 else
"000000000000" when X = 34 AND Y = 2 else
"000000000000" when X = 35 AND Y = 2 else
"000000000000" when X = 36 AND Y = 2 else
"000000000000" when X = 37 AND Y = 2 else
"000000000000" when X = 38 AND Y = 2 else
"000000000000" when X = 39 AND Y = 2 else
"000000000000" when X = 40 AND Y = 2 else
"000000000000" when X = 41 AND Y = 2 else
"000000000000" when X = 42 AND Y = 2 else
"000000000000" when X = 43 AND Y = 2 else
"000000000000" when X = 44 AND Y = 2 else
"000000000000" when X = 45 AND Y = 2 else
"000000000000" when X = 46 AND Y = 2 else
"000000000000" when X = 47 AND Y = 2 else
"000000000000" when X = 48 AND Y = 2 else
"000000000000" when X = 49 AND Y = 2 else
"000000000000" when X = 50 AND Y = 2 else
"000000000000" when X = 51 AND Y = 2 else
"000000000000" when X = 52 AND Y = 2 else
"000000000000" when X = 53 AND Y = 2 else
"000000000000" when X = 54 AND Y = 2 else
"000000000000" when X = 55 AND Y = 2 else
"000000000000" when X = 56 AND Y = 2 else
"000000000000" when X = 57 AND Y = 2 else
"000000000000" when X = 58 AND Y = 2 else
"000000000000" when X = 59 AND Y = 2 else
"000000000000" when X = 60 AND Y = 2 else
"000000000000" when X = 61 AND Y = 2 else
"000000000000" when X = 62 AND Y = 2 else
"000000000000" when X = 63 AND Y = 2 else
"000000000000" when X = 64 AND Y = 2 else
"000000000000" when X = 65 AND Y = 2 else
"000000000000" when X = 66 AND Y = 2 else
"000000000000" when X = 67 AND Y = 2 else
"000000000000" when X = 68 AND Y = 2 else
"000000000000" when X = 69 AND Y = 2 else
"000000000000" when X = 70 AND Y = 2 else
"000000000000" when X = 71 AND Y = 2 else
"000000000000" when X = 72 AND Y = 2 else
"000000000000" when X = 73 AND Y = 2 else
"000000000000" when X = 74 AND Y = 2 else
"000000000000" when X = 75 AND Y = 2 else
"000000000000" when X = 76 AND Y = 2 else
"000000000000" when X = 77 AND Y = 2 else
"000000000000" when X = 78 AND Y = 2 else
"000000000000" when X = 79 AND Y = 2 else
"111111111111" when X = 80 AND Y = 2 else
"111111111111" when X = 81 AND Y = 2 else
"111111111111" when X = 82 AND Y = 2 else
"111111111111" when X = 83 AND Y = 2 else
"111111111111" when X = 84 AND Y = 2 else
"111111111111" when X = 85 AND Y = 2 else
"111111111111" when X = 86 AND Y = 2 else
"111111111111" when X = 87 AND Y = 2 else
"111111111111" when X = 88 AND Y = 2 else
"111111111111" when X = 89 AND Y = 2 else
"111111111111" when X = 90 AND Y = 2 else
"111111111111" when X = 91 AND Y = 2 else
"111111111111" when X = 92 AND Y = 2 else
"111111111111" when X = 93 AND Y = 2 else
"111111111111" when X = 94 AND Y = 2 else
"111111111111" when X = 95 AND Y = 2 else
"111111111111" when X = 96 AND Y = 2 else
"111111111111" when X = 97 AND Y = 2 else
"111111111111" when X = 98 AND Y = 2 else
"111111111111" when X = 99 AND Y = 2 else
"111111111111" when X = 100 AND Y = 2 else
"111111111111" when X = 101 AND Y = 2 else
"111111111111" when X = 102 AND Y = 2 else
"111111111111" when X = 103 AND Y = 2 else
"111111111111" when X = 104 AND Y = 2 else
"111111111111" when X = 105 AND Y = 2 else
"111111111111" when X = 106 AND Y = 2 else
"111111111111" when X = 107 AND Y = 2 else
"111111111111" when X = 108 AND Y = 2 else
"111111111111" when X = 109 AND Y = 2 else
"111111111111" when X = 110 AND Y = 2 else
"111111111111" when X = 111 AND Y = 2 else
"111111111111" when X = 112 AND Y = 2 else
"111111111111" when X = 113 AND Y = 2 else
"111111111111" when X = 114 AND Y = 2 else
"111111111111" when X = 115 AND Y = 2 else
"111111111111" when X = 116 AND Y = 2 else
"111111111111" when X = 117 AND Y = 2 else
"111111111111" when X = 118 AND Y = 2 else
"111111111111" when X = 119 AND Y = 2 else
"111111111111" when X = 120 AND Y = 2 else
"111111111111" when X = 121 AND Y = 2 else
"111111111111" when X = 122 AND Y = 2 else
"111111111111" when X = 123 AND Y = 2 else
"111111111111" when X = 124 AND Y = 2 else
"111111111111" when X = 125 AND Y = 2 else
"111111111111" when X = 126 AND Y = 2 else
"111111111111" when X = 127 AND Y = 2 else
"111111111111" when X = 128 AND Y = 2 else
"111111111111" when X = 129 AND Y = 2 else
"111111111111" when X = 130 AND Y = 2 else
"111111111111" when X = 131 AND Y = 2 else
"111111111111" when X = 132 AND Y = 2 else
"111111111111" when X = 133 AND Y = 2 else
"111111111111" when X = 134 AND Y = 2 else
"111111111111" when X = 135 AND Y = 2 else
"111111111111" when X = 136 AND Y = 2 else
"111111111111" when X = 137 AND Y = 2 else
"111111111111" when X = 138 AND Y = 2 else
"111111111111" when X = 139 AND Y = 2 else
"000000000000" when X = 140 AND Y = 2 else
"000000000000" when X = 141 AND Y = 2 else
"000000000000" when X = 142 AND Y = 2 else
"000000000000" when X = 143 AND Y = 2 else
"000000000000" when X = 144 AND Y = 2 else
"000000000000" when X = 145 AND Y = 2 else
"000000000000" when X = 146 AND Y = 2 else
"000000000000" when X = 147 AND Y = 2 else
"000000000000" when X = 148 AND Y = 2 else
"000000000000" when X = 149 AND Y = 2 else
"000000000000" when X = 150 AND Y = 2 else
"000000000000" when X = 151 AND Y = 2 else
"000000000000" when X = 152 AND Y = 2 else
"000000000000" when X = 153 AND Y = 2 else
"000000000000" when X = 154 AND Y = 2 else
"000000000000" when X = 155 AND Y = 2 else
"000000000000" when X = 156 AND Y = 2 else
"000000000000" when X = 157 AND Y = 2 else
"000000000000" when X = 158 AND Y = 2 else
"000000000000" when X = 159 AND Y = 2 else
"000000000000" when X = 160 AND Y = 2 else
"000000000000" when X = 161 AND Y = 2 else
"000000000000" when X = 162 AND Y = 2 else
"000000000000" when X = 163 AND Y = 2 else
"000000000000" when X = 164 AND Y = 2 else
"000000000000" when X = 165 AND Y = 2 else
"000000000000" when X = 166 AND Y = 2 else
"000000000000" when X = 167 AND Y = 2 else
"000000000000" when X = 168 AND Y = 2 else
"000000000000" when X = 169 AND Y = 2 else
"000000000000" when X = 170 AND Y = 2 else
"000000000000" when X = 171 AND Y = 2 else
"000000000000" when X = 172 AND Y = 2 else
"000000000000" when X = 173 AND Y = 2 else
"000000000000" when X = 174 AND Y = 2 else
"000000000000" when X = 175 AND Y = 2 else
"000000000000" when X = 176 AND Y = 2 else
"000000000000" when X = 177 AND Y = 2 else
"000000000000" when X = 178 AND Y = 2 else
"000000000000" when X = 179 AND Y = 2 else
"000000000000" when X = 180 AND Y = 2 else
"000000000000" when X = 181 AND Y = 2 else
"000000000000" when X = 182 AND Y = 2 else
"000000000000" when X = 183 AND Y = 2 else
"000000000000" when X = 184 AND Y = 2 else
"000000000000" when X = 185 AND Y = 2 else
"000000000000" when X = 186 AND Y = 2 else
"000000000000" when X = 187 AND Y = 2 else
"000000000000" when X = 188 AND Y = 2 else
"000000000000" when X = 189 AND Y = 2 else
"000000000000" when X = 190 AND Y = 2 else
"000000000000" when X = 191 AND Y = 2 else
"000000000000" when X = 192 AND Y = 2 else
"000000000000" when X = 193 AND Y = 2 else
"000000000000" when X = 194 AND Y = 2 else
"000000000000" when X = 195 AND Y = 2 else
"000000000000" when X = 196 AND Y = 2 else
"000000000000" when X = 197 AND Y = 2 else
"000000000000" when X = 198 AND Y = 2 else
"000000000000" when X = 199 AND Y = 2 else
"000000000000" when X = 200 AND Y = 2 else
"000000000000" when X = 201 AND Y = 2 else
"000000000000" when X = 202 AND Y = 2 else
"000000000000" when X = 203 AND Y = 2 else
"000000000000" when X = 204 AND Y = 2 else
"000000000000" when X = 205 AND Y = 2 else
"000000000000" when X = 206 AND Y = 2 else
"000000000000" when X = 207 AND Y = 2 else
"000000000000" when X = 208 AND Y = 2 else
"000000000000" when X = 209 AND Y = 2 else
"000000000000" when X = 210 AND Y = 2 else
"000000000000" when X = 211 AND Y = 2 else
"000000000000" when X = 212 AND Y = 2 else
"000000000000" when X = 213 AND Y = 2 else
"000000000000" when X = 214 AND Y = 2 else
"000000000000" when X = 215 AND Y = 2 else
"000000000000" when X = 216 AND Y = 2 else
"000000000000" when X = 217 AND Y = 2 else
"000000000000" when X = 218 AND Y = 2 else
"000000000000" when X = 219 AND Y = 2 else
"000000000000" when X = 220 AND Y = 2 else
"000000000000" when X = 221 AND Y = 2 else
"000000000000" when X = 222 AND Y = 2 else
"000000000000" when X = 223 AND Y = 2 else
"000000000000" when X = 224 AND Y = 2 else
"000000000000" when X = 225 AND Y = 2 else
"000000000000" when X = 226 AND Y = 2 else
"000000000000" when X = 227 AND Y = 2 else
"000000000000" when X = 228 AND Y = 2 else
"000000000000" when X = 229 AND Y = 2 else
"000000000000" when X = 230 AND Y = 2 else
"000000000000" when X = 231 AND Y = 2 else
"000000000000" when X = 232 AND Y = 2 else
"000000000000" when X = 233 AND Y = 2 else
"000000000000" when X = 234 AND Y = 2 else
"000000000000" when X = 235 AND Y = 2 else
"000000000000" when X = 236 AND Y = 2 else
"000000000000" when X = 237 AND Y = 2 else
"000000000000" when X = 238 AND Y = 2 else
"000000000000" when X = 239 AND Y = 2 else
"000000000000" when X = 240 AND Y = 2 else
"000000000000" when X = 241 AND Y = 2 else
"000000000000" when X = 242 AND Y = 2 else
"000000000000" when X = 243 AND Y = 2 else
"000000000000" when X = 244 AND Y = 2 else
"000000000000" when X = 245 AND Y = 2 else
"000000000000" when X = 246 AND Y = 2 else
"000000000000" when X = 247 AND Y = 2 else
"000000000000" when X = 248 AND Y = 2 else
"000000000000" when X = 249 AND Y = 2 else
"000000000000" when X = 250 AND Y = 2 else
"000000000000" when X = 251 AND Y = 2 else
"000000000000" when X = 252 AND Y = 2 else
"000000000000" when X = 253 AND Y = 2 else
"000000000000" when X = 254 AND Y = 2 else
"000000000000" when X = 255 AND Y = 2 else
"000000000000" when X = 256 AND Y = 2 else
"000000000000" when X = 257 AND Y = 2 else
"000000000000" when X = 258 AND Y = 2 else
"000000000000" when X = 259 AND Y = 2 else
"000000000000" when X = 260 AND Y = 2 else
"000000000000" when X = 261 AND Y = 2 else
"000000000000" when X = 262 AND Y = 2 else
"000000000000" when X = 263 AND Y = 2 else
"000000000000" when X = 264 AND Y = 2 else
"000000000000" when X = 265 AND Y = 2 else
"000000000000" when X = 266 AND Y = 2 else
"000000000000" when X = 267 AND Y = 2 else
"000000000000" when X = 268 AND Y = 2 else
"000000000000" when X = 269 AND Y = 2 else
"000000000000" when X = 270 AND Y = 2 else
"000000000000" when X = 271 AND Y = 2 else
"000000000000" when X = 272 AND Y = 2 else
"000000000000" when X = 273 AND Y = 2 else
"000000000000" when X = 274 AND Y = 2 else
"000000000000" when X = 275 AND Y = 2 else
"000000000000" when X = 276 AND Y = 2 else
"000000000000" when X = 277 AND Y = 2 else
"000000000000" when X = 278 AND Y = 2 else
"000000000000" when X = 279 AND Y = 2 else
"000000000000" when X = 280 AND Y = 2 else
"000000000000" when X = 281 AND Y = 2 else
"000000000000" when X = 282 AND Y = 2 else
"000000000000" when X = 283 AND Y = 2 else
"000000000000" when X = 284 AND Y = 2 else
"000000000000" when X = 285 AND Y = 2 else
"000000000000" when X = 286 AND Y = 2 else
"000000000000" when X = 287 AND Y = 2 else
"000000000000" when X = 288 AND Y = 2 else
"000000000000" when X = 289 AND Y = 2 else
"000000000000" when X = 290 AND Y = 2 else
"000000000000" when X = 291 AND Y = 2 else
"000000000000" when X = 292 AND Y = 2 else
"000000000000" when X = 293 AND Y = 2 else
"000000000000" when X = 294 AND Y = 2 else
"000000000000" when X = 295 AND Y = 2 else
"000000000000" when X = 296 AND Y = 2 else
"000000000000" when X = 297 AND Y = 2 else
"000000000000" when X = 298 AND Y = 2 else
"000000000000" when X = 299 AND Y = 2 else
"000000000000" when X = 300 AND Y = 2 else
"000000000000" when X = 301 AND Y = 2 else
"000000000000" when X = 302 AND Y = 2 else
"000000000000" when X = 303 AND Y = 2 else
"000000000000" when X = 304 AND Y = 2 else
"000000000000" when X = 305 AND Y = 2 else
"000000000000" when X = 306 AND Y = 2 else
"000000000000" when X = 307 AND Y = 2 else
"000000000000" when X = 308 AND Y = 2 else
"000000000000" when X = 309 AND Y = 2 else
"000000000000" when X = 310 AND Y = 2 else
"000000000000" when X = 311 AND Y = 2 else
"000000000000" when X = 312 AND Y = 2 else
"000000000000" when X = 313 AND Y = 2 else
"000000000000" when X = 314 AND Y = 2 else
"000000000000" when X = 315 AND Y = 2 else
"000000000000" when X = 316 AND Y = 2 else
"000000000000" when X = 317 AND Y = 2 else
"000000000000" when X = 318 AND Y = 2 else
"000000000000" when X = 319 AND Y = 2 else
"000000000000" when X = 320 AND Y = 2 else
"000000000000" when X = 321 AND Y = 2 else
"000000000000" when X = 322 AND Y = 2 else
"000000000000" when X = 323 AND Y = 2 else
"000000000000" when X = 324 AND Y = 2 else
"000000000000" when X = 0 AND Y = 3 else
"000000000000" when X = 1 AND Y = 3 else
"000000000000" when X = 2 AND Y = 3 else
"000000000000" when X = 3 AND Y = 3 else
"000000000000" when X = 4 AND Y = 3 else
"000000000000" when X = 5 AND Y = 3 else
"000000000000" when X = 6 AND Y = 3 else
"000000000000" when X = 7 AND Y = 3 else
"000000000000" when X = 8 AND Y = 3 else
"000000000000" when X = 9 AND Y = 3 else
"000000000000" when X = 10 AND Y = 3 else
"000000000000" when X = 11 AND Y = 3 else
"000000000000" when X = 12 AND Y = 3 else
"000000000000" when X = 13 AND Y = 3 else
"000000000000" when X = 14 AND Y = 3 else
"000000000000" when X = 15 AND Y = 3 else
"000000000000" when X = 16 AND Y = 3 else
"000000000000" when X = 17 AND Y = 3 else
"000000000000" when X = 18 AND Y = 3 else
"000000000000" when X = 19 AND Y = 3 else
"000000000000" when X = 20 AND Y = 3 else
"000000000000" when X = 21 AND Y = 3 else
"000000000000" when X = 22 AND Y = 3 else
"000000000000" when X = 23 AND Y = 3 else
"000000000000" when X = 24 AND Y = 3 else
"000000000000" when X = 25 AND Y = 3 else
"000000000000" when X = 26 AND Y = 3 else
"000000000000" when X = 27 AND Y = 3 else
"000000000000" when X = 28 AND Y = 3 else
"000000000000" when X = 29 AND Y = 3 else
"000000000000" when X = 30 AND Y = 3 else
"000000000000" when X = 31 AND Y = 3 else
"000000000000" when X = 32 AND Y = 3 else
"000000000000" when X = 33 AND Y = 3 else
"000000000000" when X = 34 AND Y = 3 else
"000000000000" when X = 35 AND Y = 3 else
"000000000000" when X = 36 AND Y = 3 else
"000000000000" when X = 37 AND Y = 3 else
"000000000000" when X = 38 AND Y = 3 else
"000000000000" when X = 39 AND Y = 3 else
"000000000000" when X = 40 AND Y = 3 else
"000000000000" when X = 41 AND Y = 3 else
"000000000000" when X = 42 AND Y = 3 else
"000000000000" when X = 43 AND Y = 3 else
"000000000000" when X = 44 AND Y = 3 else
"000000000000" when X = 45 AND Y = 3 else
"000000000000" when X = 46 AND Y = 3 else
"000000000000" when X = 47 AND Y = 3 else
"000000000000" when X = 48 AND Y = 3 else
"000000000000" when X = 49 AND Y = 3 else
"000000000000" when X = 50 AND Y = 3 else
"000000000000" when X = 51 AND Y = 3 else
"000000000000" when X = 52 AND Y = 3 else
"000000000000" when X = 53 AND Y = 3 else
"000000000000" when X = 54 AND Y = 3 else
"000000000000" when X = 55 AND Y = 3 else
"000000000000" when X = 56 AND Y = 3 else
"000000000000" when X = 57 AND Y = 3 else
"000000000000" when X = 58 AND Y = 3 else
"000000000000" when X = 59 AND Y = 3 else
"000000000000" when X = 60 AND Y = 3 else
"000000000000" when X = 61 AND Y = 3 else
"000000000000" when X = 62 AND Y = 3 else
"000000000000" when X = 63 AND Y = 3 else
"000000000000" when X = 64 AND Y = 3 else
"000000000000" when X = 65 AND Y = 3 else
"000000000000" when X = 66 AND Y = 3 else
"000000000000" when X = 67 AND Y = 3 else
"000000000000" when X = 68 AND Y = 3 else
"000000000000" when X = 69 AND Y = 3 else
"000000000000" when X = 70 AND Y = 3 else
"000000000000" when X = 71 AND Y = 3 else
"000000000000" when X = 72 AND Y = 3 else
"000000000000" when X = 73 AND Y = 3 else
"000000000000" when X = 74 AND Y = 3 else
"000000000000" when X = 75 AND Y = 3 else
"000000000000" when X = 76 AND Y = 3 else
"000000000000" when X = 77 AND Y = 3 else
"000000000000" when X = 78 AND Y = 3 else
"000000000000" when X = 79 AND Y = 3 else
"111111111111" when X = 80 AND Y = 3 else
"111111111111" when X = 81 AND Y = 3 else
"111111111111" when X = 82 AND Y = 3 else
"111111111111" when X = 83 AND Y = 3 else
"111111111111" when X = 84 AND Y = 3 else
"111111111111" when X = 85 AND Y = 3 else
"111111111111" when X = 86 AND Y = 3 else
"111111111111" when X = 87 AND Y = 3 else
"111111111111" when X = 88 AND Y = 3 else
"111111111111" when X = 89 AND Y = 3 else
"111111111111" when X = 90 AND Y = 3 else
"111111111111" when X = 91 AND Y = 3 else
"111111111111" when X = 92 AND Y = 3 else
"111111111111" when X = 93 AND Y = 3 else
"111111111111" when X = 94 AND Y = 3 else
"111111111111" when X = 95 AND Y = 3 else
"111111111111" when X = 96 AND Y = 3 else
"111111111111" when X = 97 AND Y = 3 else
"111111111111" when X = 98 AND Y = 3 else
"111111111111" when X = 99 AND Y = 3 else
"111111111111" when X = 100 AND Y = 3 else
"111111111111" when X = 101 AND Y = 3 else
"111111111111" when X = 102 AND Y = 3 else
"111111111111" when X = 103 AND Y = 3 else
"111111111111" when X = 104 AND Y = 3 else
"111111111111" when X = 105 AND Y = 3 else
"111111111111" when X = 106 AND Y = 3 else
"111111111111" when X = 107 AND Y = 3 else
"111111111111" when X = 108 AND Y = 3 else
"111111111111" when X = 109 AND Y = 3 else
"111111111111" when X = 110 AND Y = 3 else
"111111111111" when X = 111 AND Y = 3 else
"111111111111" when X = 112 AND Y = 3 else
"111111111111" when X = 113 AND Y = 3 else
"111111111111" when X = 114 AND Y = 3 else
"111111111111" when X = 115 AND Y = 3 else
"111111111111" when X = 116 AND Y = 3 else
"111111111111" when X = 117 AND Y = 3 else
"111111111111" when X = 118 AND Y = 3 else
"111111111111" when X = 119 AND Y = 3 else
"111111111111" when X = 120 AND Y = 3 else
"111111111111" when X = 121 AND Y = 3 else
"111111111111" when X = 122 AND Y = 3 else
"111111111111" when X = 123 AND Y = 3 else
"111111111111" when X = 124 AND Y = 3 else
"111111111111" when X = 125 AND Y = 3 else
"111111111111" when X = 126 AND Y = 3 else
"111111111111" when X = 127 AND Y = 3 else
"111111111111" when X = 128 AND Y = 3 else
"111111111111" when X = 129 AND Y = 3 else
"111111111111" when X = 130 AND Y = 3 else
"111111111111" when X = 131 AND Y = 3 else
"111111111111" when X = 132 AND Y = 3 else
"111111111111" when X = 133 AND Y = 3 else
"111111111111" when X = 134 AND Y = 3 else
"111111111111" when X = 135 AND Y = 3 else
"111111111111" when X = 136 AND Y = 3 else
"111111111111" when X = 137 AND Y = 3 else
"111111111111" when X = 138 AND Y = 3 else
"111111111111" when X = 139 AND Y = 3 else
"000000000000" when X = 140 AND Y = 3 else
"000000000000" when X = 141 AND Y = 3 else
"000000000000" when X = 142 AND Y = 3 else
"000000000000" when X = 143 AND Y = 3 else
"000000000000" when X = 144 AND Y = 3 else
"000000000000" when X = 145 AND Y = 3 else
"000000000000" when X = 146 AND Y = 3 else
"000000000000" when X = 147 AND Y = 3 else
"000000000000" when X = 148 AND Y = 3 else
"000000000000" when X = 149 AND Y = 3 else
"000000000000" when X = 150 AND Y = 3 else
"000000000000" when X = 151 AND Y = 3 else
"000000000000" when X = 152 AND Y = 3 else
"000000000000" when X = 153 AND Y = 3 else
"000000000000" when X = 154 AND Y = 3 else
"000000000000" when X = 155 AND Y = 3 else
"000000000000" when X = 156 AND Y = 3 else
"000000000000" when X = 157 AND Y = 3 else
"000000000000" when X = 158 AND Y = 3 else
"000000000000" when X = 159 AND Y = 3 else
"000000000000" when X = 160 AND Y = 3 else
"000000000000" when X = 161 AND Y = 3 else
"000000000000" when X = 162 AND Y = 3 else
"000000000000" when X = 163 AND Y = 3 else
"000000000000" when X = 164 AND Y = 3 else
"000000000000" when X = 165 AND Y = 3 else
"000000000000" when X = 166 AND Y = 3 else
"000000000000" when X = 167 AND Y = 3 else
"000000000000" when X = 168 AND Y = 3 else
"000000000000" when X = 169 AND Y = 3 else
"000000000000" when X = 170 AND Y = 3 else
"000000000000" when X = 171 AND Y = 3 else
"000000000000" when X = 172 AND Y = 3 else
"000000000000" when X = 173 AND Y = 3 else
"000000000000" when X = 174 AND Y = 3 else
"000000000000" when X = 175 AND Y = 3 else
"000000000000" when X = 176 AND Y = 3 else
"000000000000" when X = 177 AND Y = 3 else
"000000000000" when X = 178 AND Y = 3 else
"000000000000" when X = 179 AND Y = 3 else
"000000000000" when X = 180 AND Y = 3 else
"000000000000" when X = 181 AND Y = 3 else
"000000000000" when X = 182 AND Y = 3 else
"000000000000" when X = 183 AND Y = 3 else
"000000000000" when X = 184 AND Y = 3 else
"000000000000" when X = 185 AND Y = 3 else
"000000000000" when X = 186 AND Y = 3 else
"000000000000" when X = 187 AND Y = 3 else
"000000000000" when X = 188 AND Y = 3 else
"000000000000" when X = 189 AND Y = 3 else
"000000000000" when X = 190 AND Y = 3 else
"000000000000" when X = 191 AND Y = 3 else
"000000000000" when X = 192 AND Y = 3 else
"000000000000" when X = 193 AND Y = 3 else
"000000000000" when X = 194 AND Y = 3 else
"000000000000" when X = 195 AND Y = 3 else
"000000000000" when X = 196 AND Y = 3 else
"000000000000" when X = 197 AND Y = 3 else
"000000000000" when X = 198 AND Y = 3 else
"000000000000" when X = 199 AND Y = 3 else
"000000000000" when X = 200 AND Y = 3 else
"000000000000" when X = 201 AND Y = 3 else
"000000000000" when X = 202 AND Y = 3 else
"000000000000" when X = 203 AND Y = 3 else
"000000000000" when X = 204 AND Y = 3 else
"000000000000" when X = 205 AND Y = 3 else
"000000000000" when X = 206 AND Y = 3 else
"000000000000" when X = 207 AND Y = 3 else
"000000000000" when X = 208 AND Y = 3 else
"000000000000" when X = 209 AND Y = 3 else
"000000000000" when X = 210 AND Y = 3 else
"000000000000" when X = 211 AND Y = 3 else
"000000000000" when X = 212 AND Y = 3 else
"000000000000" when X = 213 AND Y = 3 else
"000000000000" when X = 214 AND Y = 3 else
"000000000000" when X = 215 AND Y = 3 else
"000000000000" when X = 216 AND Y = 3 else
"000000000000" when X = 217 AND Y = 3 else
"000000000000" when X = 218 AND Y = 3 else
"000000000000" when X = 219 AND Y = 3 else
"000000000000" when X = 220 AND Y = 3 else
"000000000000" when X = 221 AND Y = 3 else
"000000000000" when X = 222 AND Y = 3 else
"000000000000" when X = 223 AND Y = 3 else
"000000000000" when X = 224 AND Y = 3 else
"000000000000" when X = 225 AND Y = 3 else
"000000000000" when X = 226 AND Y = 3 else
"000000000000" when X = 227 AND Y = 3 else
"000000000000" when X = 228 AND Y = 3 else
"000000000000" when X = 229 AND Y = 3 else
"000000000000" when X = 230 AND Y = 3 else
"000000000000" when X = 231 AND Y = 3 else
"000000000000" when X = 232 AND Y = 3 else
"000000000000" when X = 233 AND Y = 3 else
"000000000000" when X = 234 AND Y = 3 else
"000000000000" when X = 235 AND Y = 3 else
"000000000000" when X = 236 AND Y = 3 else
"000000000000" when X = 237 AND Y = 3 else
"000000000000" when X = 238 AND Y = 3 else
"000000000000" when X = 239 AND Y = 3 else
"000000000000" when X = 240 AND Y = 3 else
"000000000000" when X = 241 AND Y = 3 else
"000000000000" when X = 242 AND Y = 3 else
"000000000000" when X = 243 AND Y = 3 else
"000000000000" when X = 244 AND Y = 3 else
"000000000000" when X = 245 AND Y = 3 else
"000000000000" when X = 246 AND Y = 3 else
"000000000000" when X = 247 AND Y = 3 else
"000000000000" when X = 248 AND Y = 3 else
"000000000000" when X = 249 AND Y = 3 else
"000000000000" when X = 250 AND Y = 3 else
"000000000000" when X = 251 AND Y = 3 else
"000000000000" when X = 252 AND Y = 3 else
"000000000000" when X = 253 AND Y = 3 else
"000000000000" when X = 254 AND Y = 3 else
"000000000000" when X = 255 AND Y = 3 else
"000000000000" when X = 256 AND Y = 3 else
"000000000000" when X = 257 AND Y = 3 else
"000000000000" when X = 258 AND Y = 3 else
"000000000000" when X = 259 AND Y = 3 else
"000000000000" when X = 260 AND Y = 3 else
"000000000000" when X = 261 AND Y = 3 else
"000000000000" when X = 262 AND Y = 3 else
"000000000000" when X = 263 AND Y = 3 else
"000000000000" when X = 264 AND Y = 3 else
"000000000000" when X = 265 AND Y = 3 else
"000000000000" when X = 266 AND Y = 3 else
"000000000000" when X = 267 AND Y = 3 else
"000000000000" when X = 268 AND Y = 3 else
"000000000000" when X = 269 AND Y = 3 else
"000000000000" when X = 270 AND Y = 3 else
"000000000000" when X = 271 AND Y = 3 else
"000000000000" when X = 272 AND Y = 3 else
"000000000000" when X = 273 AND Y = 3 else
"000000000000" when X = 274 AND Y = 3 else
"000000000000" when X = 275 AND Y = 3 else
"000000000000" when X = 276 AND Y = 3 else
"000000000000" when X = 277 AND Y = 3 else
"000000000000" when X = 278 AND Y = 3 else
"000000000000" when X = 279 AND Y = 3 else
"000000000000" when X = 280 AND Y = 3 else
"000000000000" when X = 281 AND Y = 3 else
"000000000000" when X = 282 AND Y = 3 else
"000000000000" when X = 283 AND Y = 3 else
"000000000000" when X = 284 AND Y = 3 else
"000000000000" when X = 285 AND Y = 3 else
"000000000000" when X = 286 AND Y = 3 else
"000000000000" when X = 287 AND Y = 3 else
"000000000000" when X = 288 AND Y = 3 else
"000000000000" when X = 289 AND Y = 3 else
"000000000000" when X = 290 AND Y = 3 else
"000000000000" when X = 291 AND Y = 3 else
"000000000000" when X = 292 AND Y = 3 else
"000000000000" when X = 293 AND Y = 3 else
"000000000000" when X = 294 AND Y = 3 else
"000000000000" when X = 295 AND Y = 3 else
"000000000000" when X = 296 AND Y = 3 else
"000000000000" when X = 297 AND Y = 3 else
"000000000000" when X = 298 AND Y = 3 else
"000000000000" when X = 299 AND Y = 3 else
"000000000000" when X = 300 AND Y = 3 else
"000000000000" when X = 301 AND Y = 3 else
"000000000000" when X = 302 AND Y = 3 else
"000000000000" when X = 303 AND Y = 3 else
"000000000000" when X = 304 AND Y = 3 else
"000000000000" when X = 305 AND Y = 3 else
"000000000000" when X = 306 AND Y = 3 else
"000000000000" when X = 307 AND Y = 3 else
"000000000000" when X = 308 AND Y = 3 else
"000000000000" when X = 309 AND Y = 3 else
"000000000000" when X = 310 AND Y = 3 else
"000000000000" when X = 311 AND Y = 3 else
"000000000000" when X = 312 AND Y = 3 else
"000000000000" when X = 313 AND Y = 3 else
"000000000000" when X = 314 AND Y = 3 else
"000000000000" when X = 315 AND Y = 3 else
"000000000000" when X = 316 AND Y = 3 else
"000000000000" when X = 317 AND Y = 3 else
"000000000000" when X = 318 AND Y = 3 else
"000000000000" when X = 319 AND Y = 3 else
"000000000000" when X = 320 AND Y = 3 else
"000000000000" when X = 321 AND Y = 3 else
"000000000000" when X = 322 AND Y = 3 else
"000000000000" when X = 323 AND Y = 3 else
"000000000000" when X = 324 AND Y = 3 else
"000000000000" when X = 0 AND Y = 4 else
"000000000000" when X = 1 AND Y = 4 else
"000000000000" when X = 2 AND Y = 4 else
"000000000000" when X = 3 AND Y = 4 else
"000000000000" when X = 4 AND Y = 4 else
"000000000000" when X = 5 AND Y = 4 else
"000000000000" when X = 6 AND Y = 4 else
"000000000000" when X = 7 AND Y = 4 else
"000000000000" when X = 8 AND Y = 4 else
"000000000000" when X = 9 AND Y = 4 else
"000000000000" when X = 10 AND Y = 4 else
"000000000000" when X = 11 AND Y = 4 else
"000000000000" when X = 12 AND Y = 4 else
"000000000000" when X = 13 AND Y = 4 else
"000000000000" when X = 14 AND Y = 4 else
"000000000000" when X = 15 AND Y = 4 else
"000000000000" when X = 16 AND Y = 4 else
"000000000000" when X = 17 AND Y = 4 else
"000000000000" when X = 18 AND Y = 4 else
"000000000000" when X = 19 AND Y = 4 else
"000000000000" when X = 20 AND Y = 4 else
"000000000000" when X = 21 AND Y = 4 else
"000000000000" when X = 22 AND Y = 4 else
"000000000000" when X = 23 AND Y = 4 else
"000000000000" when X = 24 AND Y = 4 else
"000000000000" when X = 25 AND Y = 4 else
"000000000000" when X = 26 AND Y = 4 else
"000000000000" when X = 27 AND Y = 4 else
"000000000000" when X = 28 AND Y = 4 else
"000000000000" when X = 29 AND Y = 4 else
"000000000000" when X = 30 AND Y = 4 else
"000000000000" when X = 31 AND Y = 4 else
"000000000000" when X = 32 AND Y = 4 else
"000000000000" when X = 33 AND Y = 4 else
"000000000000" when X = 34 AND Y = 4 else
"000000000000" when X = 35 AND Y = 4 else
"000000000000" when X = 36 AND Y = 4 else
"000000000000" when X = 37 AND Y = 4 else
"000000000000" when X = 38 AND Y = 4 else
"000000000000" when X = 39 AND Y = 4 else
"000000000000" when X = 40 AND Y = 4 else
"000000000000" when X = 41 AND Y = 4 else
"000000000000" when X = 42 AND Y = 4 else
"000000000000" when X = 43 AND Y = 4 else
"000000000000" when X = 44 AND Y = 4 else
"000000000000" when X = 45 AND Y = 4 else
"000000000000" when X = 46 AND Y = 4 else
"000000000000" when X = 47 AND Y = 4 else
"000000000000" when X = 48 AND Y = 4 else
"000000000000" when X = 49 AND Y = 4 else
"000000000000" when X = 50 AND Y = 4 else
"000000000000" when X = 51 AND Y = 4 else
"000000000000" when X = 52 AND Y = 4 else
"000000000000" when X = 53 AND Y = 4 else
"000000000000" when X = 54 AND Y = 4 else
"000000000000" when X = 55 AND Y = 4 else
"000000000000" when X = 56 AND Y = 4 else
"000000000000" when X = 57 AND Y = 4 else
"000000000000" when X = 58 AND Y = 4 else
"000000000000" when X = 59 AND Y = 4 else
"000000000000" when X = 60 AND Y = 4 else
"000000000000" when X = 61 AND Y = 4 else
"000000000000" when X = 62 AND Y = 4 else
"000000000000" when X = 63 AND Y = 4 else
"000000000000" when X = 64 AND Y = 4 else
"000000000000" when X = 65 AND Y = 4 else
"000000000000" when X = 66 AND Y = 4 else
"000000000000" when X = 67 AND Y = 4 else
"000000000000" when X = 68 AND Y = 4 else
"000000000000" when X = 69 AND Y = 4 else
"000000000000" when X = 70 AND Y = 4 else
"000000000000" when X = 71 AND Y = 4 else
"000000000000" when X = 72 AND Y = 4 else
"000000000000" when X = 73 AND Y = 4 else
"000000000000" when X = 74 AND Y = 4 else
"000000000000" when X = 75 AND Y = 4 else
"000000000000" when X = 76 AND Y = 4 else
"000000000000" when X = 77 AND Y = 4 else
"000000000000" when X = 78 AND Y = 4 else
"000000000000" when X = 79 AND Y = 4 else
"111111111111" when X = 80 AND Y = 4 else
"111111111111" when X = 81 AND Y = 4 else
"111111111111" when X = 82 AND Y = 4 else
"111111111111" when X = 83 AND Y = 4 else
"111111111111" when X = 84 AND Y = 4 else
"111111111111" when X = 85 AND Y = 4 else
"111111111111" when X = 86 AND Y = 4 else
"111111111111" when X = 87 AND Y = 4 else
"111111111111" when X = 88 AND Y = 4 else
"111111111111" when X = 89 AND Y = 4 else
"111111111111" when X = 90 AND Y = 4 else
"111111111111" when X = 91 AND Y = 4 else
"111111111111" when X = 92 AND Y = 4 else
"111111111111" when X = 93 AND Y = 4 else
"111111111111" when X = 94 AND Y = 4 else
"111111111111" when X = 95 AND Y = 4 else
"111111111111" when X = 96 AND Y = 4 else
"111111111111" when X = 97 AND Y = 4 else
"111111111111" when X = 98 AND Y = 4 else
"111111111111" when X = 99 AND Y = 4 else
"111111111111" when X = 100 AND Y = 4 else
"111111111111" when X = 101 AND Y = 4 else
"111111111111" when X = 102 AND Y = 4 else
"111111111111" when X = 103 AND Y = 4 else
"111111111111" when X = 104 AND Y = 4 else
"111111111111" when X = 105 AND Y = 4 else
"111111111111" when X = 106 AND Y = 4 else
"111111111111" when X = 107 AND Y = 4 else
"111111111111" when X = 108 AND Y = 4 else
"111111111111" when X = 109 AND Y = 4 else
"111111111111" when X = 110 AND Y = 4 else
"111111111111" when X = 111 AND Y = 4 else
"111111111111" when X = 112 AND Y = 4 else
"111111111111" when X = 113 AND Y = 4 else
"111111111111" when X = 114 AND Y = 4 else
"111111111111" when X = 115 AND Y = 4 else
"111111111111" when X = 116 AND Y = 4 else
"111111111111" when X = 117 AND Y = 4 else
"111111111111" when X = 118 AND Y = 4 else
"111111111111" when X = 119 AND Y = 4 else
"111111111111" when X = 120 AND Y = 4 else
"111111111111" when X = 121 AND Y = 4 else
"111111111111" when X = 122 AND Y = 4 else
"111111111111" when X = 123 AND Y = 4 else
"111111111111" when X = 124 AND Y = 4 else
"111111111111" when X = 125 AND Y = 4 else
"111111111111" when X = 126 AND Y = 4 else
"111111111111" when X = 127 AND Y = 4 else
"111111111111" when X = 128 AND Y = 4 else
"111111111111" when X = 129 AND Y = 4 else
"111111111111" when X = 130 AND Y = 4 else
"111111111111" when X = 131 AND Y = 4 else
"111111111111" when X = 132 AND Y = 4 else
"111111111111" when X = 133 AND Y = 4 else
"111111111111" when X = 134 AND Y = 4 else
"111111111111" when X = 135 AND Y = 4 else
"111111111111" when X = 136 AND Y = 4 else
"111111111111" when X = 137 AND Y = 4 else
"111111111111" when X = 138 AND Y = 4 else
"111111111111" when X = 139 AND Y = 4 else
"000000000000" when X = 140 AND Y = 4 else
"000000000000" when X = 141 AND Y = 4 else
"000000000000" when X = 142 AND Y = 4 else
"000000000000" when X = 143 AND Y = 4 else
"000000000000" when X = 144 AND Y = 4 else
"000000000000" when X = 145 AND Y = 4 else
"000000000000" when X = 146 AND Y = 4 else
"000000000000" when X = 147 AND Y = 4 else
"000000000000" when X = 148 AND Y = 4 else
"000000000000" when X = 149 AND Y = 4 else
"000000000000" when X = 150 AND Y = 4 else
"000000000000" when X = 151 AND Y = 4 else
"000000000000" when X = 152 AND Y = 4 else
"000000000000" when X = 153 AND Y = 4 else
"000000000000" when X = 154 AND Y = 4 else
"000000000000" when X = 155 AND Y = 4 else
"000000000000" when X = 156 AND Y = 4 else
"000000000000" when X = 157 AND Y = 4 else
"000000000000" when X = 158 AND Y = 4 else
"000000000000" when X = 159 AND Y = 4 else
"000000000000" when X = 160 AND Y = 4 else
"000000000000" when X = 161 AND Y = 4 else
"000000000000" when X = 162 AND Y = 4 else
"000000000000" when X = 163 AND Y = 4 else
"000000000000" when X = 164 AND Y = 4 else
"000000000000" when X = 165 AND Y = 4 else
"000000000000" when X = 166 AND Y = 4 else
"000000000000" when X = 167 AND Y = 4 else
"000000000000" when X = 168 AND Y = 4 else
"000000000000" when X = 169 AND Y = 4 else
"000000000000" when X = 170 AND Y = 4 else
"000000000000" when X = 171 AND Y = 4 else
"000000000000" when X = 172 AND Y = 4 else
"000000000000" when X = 173 AND Y = 4 else
"000000000000" when X = 174 AND Y = 4 else
"000000000000" when X = 175 AND Y = 4 else
"000000000000" when X = 176 AND Y = 4 else
"000000000000" when X = 177 AND Y = 4 else
"000000000000" when X = 178 AND Y = 4 else
"000000000000" when X = 179 AND Y = 4 else
"000000000000" when X = 180 AND Y = 4 else
"000000000000" when X = 181 AND Y = 4 else
"000000000000" when X = 182 AND Y = 4 else
"000000000000" when X = 183 AND Y = 4 else
"000000000000" when X = 184 AND Y = 4 else
"000000000000" when X = 185 AND Y = 4 else
"000000000000" when X = 186 AND Y = 4 else
"000000000000" when X = 187 AND Y = 4 else
"000000000000" when X = 188 AND Y = 4 else
"000000000000" when X = 189 AND Y = 4 else
"000000000000" when X = 190 AND Y = 4 else
"000000000000" when X = 191 AND Y = 4 else
"000000000000" when X = 192 AND Y = 4 else
"000000000000" when X = 193 AND Y = 4 else
"000000000000" when X = 194 AND Y = 4 else
"000000000000" when X = 195 AND Y = 4 else
"000000000000" when X = 196 AND Y = 4 else
"000000000000" when X = 197 AND Y = 4 else
"000000000000" when X = 198 AND Y = 4 else
"000000000000" when X = 199 AND Y = 4 else
"000000000000" when X = 200 AND Y = 4 else
"000000000000" when X = 201 AND Y = 4 else
"000000000000" when X = 202 AND Y = 4 else
"000000000000" when X = 203 AND Y = 4 else
"000000000000" when X = 204 AND Y = 4 else
"000000000000" when X = 205 AND Y = 4 else
"000000000000" when X = 206 AND Y = 4 else
"000000000000" when X = 207 AND Y = 4 else
"000000000000" when X = 208 AND Y = 4 else
"000000000000" when X = 209 AND Y = 4 else
"000000000000" when X = 210 AND Y = 4 else
"000000000000" when X = 211 AND Y = 4 else
"000000000000" when X = 212 AND Y = 4 else
"000000000000" when X = 213 AND Y = 4 else
"000000000000" when X = 214 AND Y = 4 else
"000000000000" when X = 215 AND Y = 4 else
"000000000000" when X = 216 AND Y = 4 else
"000000000000" when X = 217 AND Y = 4 else
"000000000000" when X = 218 AND Y = 4 else
"000000000000" when X = 219 AND Y = 4 else
"000000000000" when X = 220 AND Y = 4 else
"000000000000" when X = 221 AND Y = 4 else
"000000000000" when X = 222 AND Y = 4 else
"000000000000" when X = 223 AND Y = 4 else
"000000000000" when X = 224 AND Y = 4 else
"000000000000" when X = 225 AND Y = 4 else
"000000000000" when X = 226 AND Y = 4 else
"000000000000" when X = 227 AND Y = 4 else
"000000000000" when X = 228 AND Y = 4 else
"000000000000" when X = 229 AND Y = 4 else
"000000000000" when X = 230 AND Y = 4 else
"000000000000" when X = 231 AND Y = 4 else
"000000000000" when X = 232 AND Y = 4 else
"000000000000" when X = 233 AND Y = 4 else
"000000000000" when X = 234 AND Y = 4 else
"000000000000" when X = 235 AND Y = 4 else
"000000000000" when X = 236 AND Y = 4 else
"000000000000" when X = 237 AND Y = 4 else
"000000000000" when X = 238 AND Y = 4 else
"000000000000" when X = 239 AND Y = 4 else
"000000000000" when X = 240 AND Y = 4 else
"000000000000" when X = 241 AND Y = 4 else
"000000000000" when X = 242 AND Y = 4 else
"000000000000" when X = 243 AND Y = 4 else
"000000000000" when X = 244 AND Y = 4 else
"000000000000" when X = 245 AND Y = 4 else
"000000000000" when X = 246 AND Y = 4 else
"000000000000" when X = 247 AND Y = 4 else
"000000000000" when X = 248 AND Y = 4 else
"000000000000" when X = 249 AND Y = 4 else
"000000000000" when X = 250 AND Y = 4 else
"000000000000" when X = 251 AND Y = 4 else
"000000000000" when X = 252 AND Y = 4 else
"000000000000" when X = 253 AND Y = 4 else
"000000000000" when X = 254 AND Y = 4 else
"000000000000" when X = 255 AND Y = 4 else
"000000000000" when X = 256 AND Y = 4 else
"000000000000" when X = 257 AND Y = 4 else
"000000000000" when X = 258 AND Y = 4 else
"000000000000" when X = 259 AND Y = 4 else
"000000000000" when X = 260 AND Y = 4 else
"000000000000" when X = 261 AND Y = 4 else
"000000000000" when X = 262 AND Y = 4 else
"000000000000" when X = 263 AND Y = 4 else
"000000000000" when X = 264 AND Y = 4 else
"000000000000" when X = 265 AND Y = 4 else
"000000000000" when X = 266 AND Y = 4 else
"000000000000" when X = 267 AND Y = 4 else
"000000000000" when X = 268 AND Y = 4 else
"000000000000" when X = 269 AND Y = 4 else
"000000000000" when X = 270 AND Y = 4 else
"000000000000" when X = 271 AND Y = 4 else
"000000000000" when X = 272 AND Y = 4 else
"000000000000" when X = 273 AND Y = 4 else
"000000000000" when X = 274 AND Y = 4 else
"000000000000" when X = 275 AND Y = 4 else
"000000000000" when X = 276 AND Y = 4 else
"000000000000" when X = 277 AND Y = 4 else
"000000000000" when X = 278 AND Y = 4 else
"000000000000" when X = 279 AND Y = 4 else
"000000000000" when X = 280 AND Y = 4 else
"000000000000" when X = 281 AND Y = 4 else
"000000000000" when X = 282 AND Y = 4 else
"000000000000" when X = 283 AND Y = 4 else
"000000000000" when X = 284 AND Y = 4 else
"000000000000" when X = 285 AND Y = 4 else
"000000000000" when X = 286 AND Y = 4 else
"000000000000" when X = 287 AND Y = 4 else
"000000000000" when X = 288 AND Y = 4 else
"000000000000" when X = 289 AND Y = 4 else
"000000000000" when X = 290 AND Y = 4 else
"000000000000" when X = 291 AND Y = 4 else
"000000000000" when X = 292 AND Y = 4 else
"000000000000" when X = 293 AND Y = 4 else
"000000000000" when X = 294 AND Y = 4 else
"000000000000" when X = 295 AND Y = 4 else
"000000000000" when X = 296 AND Y = 4 else
"000000000000" when X = 297 AND Y = 4 else
"000000000000" when X = 298 AND Y = 4 else
"000000000000" when X = 299 AND Y = 4 else
"000000000000" when X = 300 AND Y = 4 else
"000000000000" when X = 301 AND Y = 4 else
"000000000000" when X = 302 AND Y = 4 else
"000000000000" when X = 303 AND Y = 4 else
"000000000000" when X = 304 AND Y = 4 else
"000000000000" when X = 305 AND Y = 4 else
"000000000000" when X = 306 AND Y = 4 else
"000000000000" when X = 307 AND Y = 4 else
"000000000000" when X = 308 AND Y = 4 else
"000000000000" when X = 309 AND Y = 4 else
"000000000000" when X = 310 AND Y = 4 else
"000000000000" when X = 311 AND Y = 4 else
"000000000000" when X = 312 AND Y = 4 else
"000000000000" when X = 313 AND Y = 4 else
"000000000000" when X = 314 AND Y = 4 else
"000000000000" when X = 315 AND Y = 4 else
"000000000000" when X = 316 AND Y = 4 else
"000000000000" when X = 317 AND Y = 4 else
"000000000000" when X = 318 AND Y = 4 else
"000000000000" when X = 319 AND Y = 4 else
"000000000000" when X = 320 AND Y = 4 else
"000000000000" when X = 321 AND Y = 4 else
"000000000000" when X = 322 AND Y = 4 else
"000000000000" when X = 323 AND Y = 4 else
"000000000000" when X = 324 AND Y = 4 else
"000000000000" when X = 0 AND Y = 5 else
"000000000000" when X = 1 AND Y = 5 else
"000000000000" when X = 2 AND Y = 5 else
"000000000000" when X = 3 AND Y = 5 else
"000000000000" when X = 4 AND Y = 5 else
"000000000000" when X = 5 AND Y = 5 else
"000000000000" when X = 6 AND Y = 5 else
"000000000000" when X = 7 AND Y = 5 else
"000000000000" when X = 8 AND Y = 5 else
"000000000000" when X = 9 AND Y = 5 else
"000000000000" when X = 10 AND Y = 5 else
"000000000000" when X = 11 AND Y = 5 else
"000000000000" when X = 12 AND Y = 5 else
"000000000000" when X = 13 AND Y = 5 else
"000000000000" when X = 14 AND Y = 5 else
"000000000000" when X = 15 AND Y = 5 else
"000000000000" when X = 16 AND Y = 5 else
"000000000000" when X = 17 AND Y = 5 else
"000000000000" when X = 18 AND Y = 5 else
"000000000000" when X = 19 AND Y = 5 else
"000000000000" when X = 20 AND Y = 5 else
"000000000000" when X = 21 AND Y = 5 else
"000000000000" when X = 22 AND Y = 5 else
"000000000000" when X = 23 AND Y = 5 else
"000000000000" when X = 24 AND Y = 5 else
"000000000000" when X = 25 AND Y = 5 else
"000000000000" when X = 26 AND Y = 5 else
"000000000000" when X = 27 AND Y = 5 else
"000000000000" when X = 28 AND Y = 5 else
"000000000000" when X = 29 AND Y = 5 else
"000000000000" when X = 30 AND Y = 5 else
"000000000000" when X = 31 AND Y = 5 else
"000000000000" when X = 32 AND Y = 5 else
"000000000000" when X = 33 AND Y = 5 else
"000000000000" when X = 34 AND Y = 5 else
"000000000000" when X = 35 AND Y = 5 else
"000000000000" when X = 36 AND Y = 5 else
"000000000000" when X = 37 AND Y = 5 else
"000000000000" when X = 38 AND Y = 5 else
"000000000000" when X = 39 AND Y = 5 else
"110111011111" when X = 40 AND Y = 5 else
"110111011111" when X = 41 AND Y = 5 else
"110111011111" when X = 42 AND Y = 5 else
"110111011111" when X = 43 AND Y = 5 else
"110111011111" when X = 44 AND Y = 5 else
"110111011111" when X = 45 AND Y = 5 else
"110111011111" when X = 46 AND Y = 5 else
"110111011111" when X = 47 AND Y = 5 else
"110111011111" when X = 48 AND Y = 5 else
"110111011111" when X = 49 AND Y = 5 else
"110111011111" when X = 50 AND Y = 5 else
"110111011111" when X = 51 AND Y = 5 else
"110111011111" when X = 52 AND Y = 5 else
"110111011111" when X = 53 AND Y = 5 else
"110111011111" when X = 54 AND Y = 5 else
"110111011111" when X = 55 AND Y = 5 else
"110111011111" when X = 56 AND Y = 5 else
"110111011111" when X = 57 AND Y = 5 else
"110111011111" when X = 58 AND Y = 5 else
"110111011111" when X = 59 AND Y = 5 else
"110111011111" when X = 60 AND Y = 5 else
"110111011111" when X = 61 AND Y = 5 else
"110111011111" when X = 62 AND Y = 5 else
"110111011111" when X = 63 AND Y = 5 else
"110111011111" when X = 64 AND Y = 5 else
"110111011111" when X = 65 AND Y = 5 else
"110111011111" when X = 66 AND Y = 5 else
"110111011111" when X = 67 AND Y = 5 else
"110111011111" when X = 68 AND Y = 5 else
"110111011111" when X = 69 AND Y = 5 else
"110111011111" when X = 70 AND Y = 5 else
"110111011111" when X = 71 AND Y = 5 else
"110111011111" when X = 72 AND Y = 5 else
"110111011111" when X = 73 AND Y = 5 else
"110111011111" when X = 74 AND Y = 5 else
"111111111111" when X = 75 AND Y = 5 else
"111111111111" when X = 76 AND Y = 5 else
"111111111111" when X = 77 AND Y = 5 else
"111111111111" when X = 78 AND Y = 5 else
"111111111111" when X = 79 AND Y = 5 else
"111111111111" when X = 80 AND Y = 5 else
"111111111111" when X = 81 AND Y = 5 else
"111111111111" when X = 82 AND Y = 5 else
"111111111111" when X = 83 AND Y = 5 else
"111111111111" when X = 84 AND Y = 5 else
"111111111111" when X = 85 AND Y = 5 else
"111111111111" when X = 86 AND Y = 5 else
"111111111111" when X = 87 AND Y = 5 else
"111111111111" when X = 88 AND Y = 5 else
"111111111111" when X = 89 AND Y = 5 else
"111111111111" when X = 90 AND Y = 5 else
"111111111111" when X = 91 AND Y = 5 else
"111111111111" when X = 92 AND Y = 5 else
"111111111111" when X = 93 AND Y = 5 else
"111111111111" when X = 94 AND Y = 5 else
"111111111111" when X = 95 AND Y = 5 else
"111111111111" when X = 96 AND Y = 5 else
"111111111111" when X = 97 AND Y = 5 else
"111111111111" when X = 98 AND Y = 5 else
"111111111111" when X = 99 AND Y = 5 else
"111111111111" when X = 100 AND Y = 5 else
"111111111111" when X = 101 AND Y = 5 else
"111111111111" when X = 102 AND Y = 5 else
"111111111111" when X = 103 AND Y = 5 else
"111111111111" when X = 104 AND Y = 5 else
"111111111111" when X = 105 AND Y = 5 else
"111111111111" when X = 106 AND Y = 5 else
"111111111111" when X = 107 AND Y = 5 else
"111111111111" when X = 108 AND Y = 5 else
"111111111111" when X = 109 AND Y = 5 else
"111111111111" when X = 110 AND Y = 5 else
"111111111111" when X = 111 AND Y = 5 else
"111111111111" when X = 112 AND Y = 5 else
"111111111111" when X = 113 AND Y = 5 else
"111111111111" when X = 114 AND Y = 5 else
"111111111111" when X = 115 AND Y = 5 else
"111111111111" when X = 116 AND Y = 5 else
"111111111111" when X = 117 AND Y = 5 else
"111111111111" when X = 118 AND Y = 5 else
"111111111111" when X = 119 AND Y = 5 else
"111111111111" when X = 120 AND Y = 5 else
"111111111111" when X = 121 AND Y = 5 else
"111111111111" when X = 122 AND Y = 5 else
"111111111111" when X = 123 AND Y = 5 else
"111111111111" when X = 124 AND Y = 5 else
"111111111111" when X = 125 AND Y = 5 else
"111111111111" when X = 126 AND Y = 5 else
"111111111111" when X = 127 AND Y = 5 else
"111111111111" when X = 128 AND Y = 5 else
"111111111111" when X = 129 AND Y = 5 else
"111111111111" when X = 130 AND Y = 5 else
"111111111111" when X = 131 AND Y = 5 else
"111111111111" when X = 132 AND Y = 5 else
"111111111111" when X = 133 AND Y = 5 else
"111111111111" when X = 134 AND Y = 5 else
"111111111111" when X = 135 AND Y = 5 else
"111111111111" when X = 136 AND Y = 5 else
"111111111111" when X = 137 AND Y = 5 else
"111111111111" when X = 138 AND Y = 5 else
"111111111111" when X = 139 AND Y = 5 else
"111111111111" when X = 140 AND Y = 5 else
"111111111111" when X = 141 AND Y = 5 else
"111111111111" when X = 142 AND Y = 5 else
"111111111111" when X = 143 AND Y = 5 else
"111111111111" when X = 144 AND Y = 5 else
"000000000000" when X = 145 AND Y = 5 else
"000000000000" when X = 146 AND Y = 5 else
"000000000000" when X = 147 AND Y = 5 else
"000000000000" when X = 148 AND Y = 5 else
"000000000000" when X = 149 AND Y = 5 else
"000000000000" when X = 150 AND Y = 5 else
"000000000000" when X = 151 AND Y = 5 else
"000000000000" when X = 152 AND Y = 5 else
"000000000000" when X = 153 AND Y = 5 else
"000000000000" when X = 154 AND Y = 5 else
"000000000000" when X = 155 AND Y = 5 else
"000000000000" when X = 156 AND Y = 5 else
"000000000000" when X = 157 AND Y = 5 else
"000000000000" when X = 158 AND Y = 5 else
"000000000000" when X = 159 AND Y = 5 else
"000000000000" when X = 160 AND Y = 5 else
"000000000000" when X = 161 AND Y = 5 else
"000000000000" when X = 162 AND Y = 5 else
"000000000000" when X = 163 AND Y = 5 else
"000000000000" when X = 164 AND Y = 5 else
"000000000000" when X = 165 AND Y = 5 else
"000000000000" when X = 166 AND Y = 5 else
"000000000000" when X = 167 AND Y = 5 else
"000000000000" when X = 168 AND Y = 5 else
"000000000000" when X = 169 AND Y = 5 else
"000000000000" when X = 170 AND Y = 5 else
"000000000000" when X = 171 AND Y = 5 else
"000000000000" when X = 172 AND Y = 5 else
"000000000000" when X = 173 AND Y = 5 else
"000000000000" when X = 174 AND Y = 5 else
"000000000000" when X = 175 AND Y = 5 else
"000000000000" when X = 176 AND Y = 5 else
"000000000000" when X = 177 AND Y = 5 else
"000000000000" when X = 178 AND Y = 5 else
"000000000000" when X = 179 AND Y = 5 else
"000000000000" when X = 180 AND Y = 5 else
"000000000000" when X = 181 AND Y = 5 else
"000000000000" when X = 182 AND Y = 5 else
"000000000000" when X = 183 AND Y = 5 else
"000000000000" when X = 184 AND Y = 5 else
"000000000000" when X = 185 AND Y = 5 else
"000000000000" when X = 186 AND Y = 5 else
"000000000000" when X = 187 AND Y = 5 else
"000000000000" when X = 188 AND Y = 5 else
"000000000000" when X = 189 AND Y = 5 else
"000000000000" when X = 190 AND Y = 5 else
"000000000000" when X = 191 AND Y = 5 else
"000000000000" when X = 192 AND Y = 5 else
"000000000000" when X = 193 AND Y = 5 else
"000000000000" when X = 194 AND Y = 5 else
"000000000000" when X = 195 AND Y = 5 else
"000000000000" when X = 196 AND Y = 5 else
"000000000000" when X = 197 AND Y = 5 else
"000000000000" when X = 198 AND Y = 5 else
"000000000000" when X = 199 AND Y = 5 else
"000000000000" when X = 200 AND Y = 5 else
"000000000000" when X = 201 AND Y = 5 else
"000000000000" when X = 202 AND Y = 5 else
"000000000000" when X = 203 AND Y = 5 else
"000000000000" when X = 204 AND Y = 5 else
"000000000000" when X = 205 AND Y = 5 else
"000000000000" when X = 206 AND Y = 5 else
"000000000000" when X = 207 AND Y = 5 else
"000000000000" when X = 208 AND Y = 5 else
"000000000000" when X = 209 AND Y = 5 else
"000000000000" when X = 210 AND Y = 5 else
"000000000000" when X = 211 AND Y = 5 else
"000000000000" when X = 212 AND Y = 5 else
"000000000000" when X = 213 AND Y = 5 else
"000000000000" when X = 214 AND Y = 5 else
"000000000000" when X = 215 AND Y = 5 else
"000000000000" when X = 216 AND Y = 5 else
"000000000000" when X = 217 AND Y = 5 else
"000000000000" when X = 218 AND Y = 5 else
"000000000000" when X = 219 AND Y = 5 else
"000000000000" when X = 220 AND Y = 5 else
"000000000000" when X = 221 AND Y = 5 else
"000000000000" when X = 222 AND Y = 5 else
"000000000000" when X = 223 AND Y = 5 else
"000000000000" when X = 224 AND Y = 5 else
"000000000000" when X = 225 AND Y = 5 else
"000000000000" when X = 226 AND Y = 5 else
"000000000000" when X = 227 AND Y = 5 else
"000000000000" when X = 228 AND Y = 5 else
"000000000000" when X = 229 AND Y = 5 else
"000000000000" when X = 230 AND Y = 5 else
"000000000000" when X = 231 AND Y = 5 else
"000000000000" when X = 232 AND Y = 5 else
"000000000000" when X = 233 AND Y = 5 else
"000000000000" when X = 234 AND Y = 5 else
"000000000000" when X = 235 AND Y = 5 else
"000000000000" when X = 236 AND Y = 5 else
"000000000000" when X = 237 AND Y = 5 else
"000000000000" when X = 238 AND Y = 5 else
"000000000000" when X = 239 AND Y = 5 else
"000000000000" when X = 240 AND Y = 5 else
"000000000000" when X = 241 AND Y = 5 else
"000000000000" when X = 242 AND Y = 5 else
"000000000000" when X = 243 AND Y = 5 else
"000000000000" when X = 244 AND Y = 5 else
"000000000000" when X = 245 AND Y = 5 else
"000000000000" when X = 246 AND Y = 5 else
"000000000000" when X = 247 AND Y = 5 else
"000000000000" when X = 248 AND Y = 5 else
"000000000000" when X = 249 AND Y = 5 else
"000000000000" when X = 250 AND Y = 5 else
"000000000000" when X = 251 AND Y = 5 else
"000000000000" when X = 252 AND Y = 5 else
"000000000000" when X = 253 AND Y = 5 else
"000000000000" when X = 254 AND Y = 5 else
"000000000000" when X = 255 AND Y = 5 else
"000000000000" when X = 256 AND Y = 5 else
"000000000000" when X = 257 AND Y = 5 else
"000000000000" when X = 258 AND Y = 5 else
"000000000000" when X = 259 AND Y = 5 else
"000000000000" when X = 260 AND Y = 5 else
"000000000000" when X = 261 AND Y = 5 else
"000000000000" when X = 262 AND Y = 5 else
"000000000000" when X = 263 AND Y = 5 else
"000000000000" when X = 264 AND Y = 5 else
"000000000000" when X = 265 AND Y = 5 else
"000000000000" when X = 266 AND Y = 5 else
"000000000000" when X = 267 AND Y = 5 else
"000000000000" when X = 268 AND Y = 5 else
"000000000000" when X = 269 AND Y = 5 else
"000000000000" when X = 270 AND Y = 5 else
"000000000000" when X = 271 AND Y = 5 else
"000000000000" when X = 272 AND Y = 5 else
"000000000000" when X = 273 AND Y = 5 else
"000000000000" when X = 274 AND Y = 5 else
"000000000000" when X = 275 AND Y = 5 else
"000000000000" when X = 276 AND Y = 5 else
"000000000000" when X = 277 AND Y = 5 else
"000000000000" when X = 278 AND Y = 5 else
"000000000000" when X = 279 AND Y = 5 else
"000000000000" when X = 280 AND Y = 5 else
"000000000000" when X = 281 AND Y = 5 else
"000000000000" when X = 282 AND Y = 5 else
"000000000000" when X = 283 AND Y = 5 else
"000000000000" when X = 284 AND Y = 5 else
"000000000000" when X = 285 AND Y = 5 else
"000000000000" when X = 286 AND Y = 5 else
"000000000000" when X = 287 AND Y = 5 else
"000000000000" when X = 288 AND Y = 5 else
"000000000000" when X = 289 AND Y = 5 else
"000000000000" when X = 290 AND Y = 5 else
"000000000000" when X = 291 AND Y = 5 else
"000000000000" when X = 292 AND Y = 5 else
"000000000000" when X = 293 AND Y = 5 else
"000000000000" when X = 294 AND Y = 5 else
"000000000000" when X = 295 AND Y = 5 else
"000000000000" when X = 296 AND Y = 5 else
"000000000000" when X = 297 AND Y = 5 else
"000000000000" when X = 298 AND Y = 5 else
"000000000000" when X = 299 AND Y = 5 else
"000000000000" when X = 300 AND Y = 5 else
"000000000000" when X = 301 AND Y = 5 else
"000000000000" when X = 302 AND Y = 5 else
"000000000000" when X = 303 AND Y = 5 else
"000000000000" when X = 304 AND Y = 5 else
"000000000000" when X = 305 AND Y = 5 else
"000000000000" when X = 306 AND Y = 5 else
"000000000000" when X = 307 AND Y = 5 else
"000000000000" when X = 308 AND Y = 5 else
"000000000000" when X = 309 AND Y = 5 else
"000000000000" when X = 310 AND Y = 5 else
"000000000000" when X = 311 AND Y = 5 else
"000000000000" when X = 312 AND Y = 5 else
"000000000000" when X = 313 AND Y = 5 else
"000000000000" when X = 314 AND Y = 5 else
"000000000000" when X = 315 AND Y = 5 else
"000000000000" when X = 316 AND Y = 5 else
"000000000000" when X = 317 AND Y = 5 else
"000000000000" when X = 318 AND Y = 5 else
"000000000000" when X = 319 AND Y = 5 else
"000000000000" when X = 320 AND Y = 5 else
"000000000000" when X = 321 AND Y = 5 else
"000000000000" when X = 322 AND Y = 5 else
"000000000000" when X = 323 AND Y = 5 else
"000000000000" when X = 324 AND Y = 5 else
"000000000000" when X = 0 AND Y = 6 else
"000000000000" when X = 1 AND Y = 6 else
"000000000000" when X = 2 AND Y = 6 else
"000000000000" when X = 3 AND Y = 6 else
"000000000000" when X = 4 AND Y = 6 else
"000000000000" when X = 5 AND Y = 6 else
"000000000000" when X = 6 AND Y = 6 else
"000000000000" when X = 7 AND Y = 6 else
"000000000000" when X = 8 AND Y = 6 else
"000000000000" when X = 9 AND Y = 6 else
"000000000000" when X = 10 AND Y = 6 else
"000000000000" when X = 11 AND Y = 6 else
"000000000000" when X = 12 AND Y = 6 else
"000000000000" when X = 13 AND Y = 6 else
"000000000000" when X = 14 AND Y = 6 else
"000000000000" when X = 15 AND Y = 6 else
"000000000000" when X = 16 AND Y = 6 else
"000000000000" when X = 17 AND Y = 6 else
"000000000000" when X = 18 AND Y = 6 else
"000000000000" when X = 19 AND Y = 6 else
"000000000000" when X = 20 AND Y = 6 else
"000000000000" when X = 21 AND Y = 6 else
"000000000000" when X = 22 AND Y = 6 else
"000000000000" when X = 23 AND Y = 6 else
"000000000000" when X = 24 AND Y = 6 else
"000000000000" when X = 25 AND Y = 6 else
"000000000000" when X = 26 AND Y = 6 else
"000000000000" when X = 27 AND Y = 6 else
"000000000000" when X = 28 AND Y = 6 else
"000000000000" when X = 29 AND Y = 6 else
"000000000000" when X = 30 AND Y = 6 else
"000000000000" when X = 31 AND Y = 6 else
"000000000000" when X = 32 AND Y = 6 else
"000000000000" when X = 33 AND Y = 6 else
"000000000000" when X = 34 AND Y = 6 else
"000000000000" when X = 35 AND Y = 6 else
"000000000000" when X = 36 AND Y = 6 else
"000000000000" when X = 37 AND Y = 6 else
"000000000000" when X = 38 AND Y = 6 else
"000000000000" when X = 39 AND Y = 6 else
"110111011111" when X = 40 AND Y = 6 else
"110111011111" when X = 41 AND Y = 6 else
"110111011111" when X = 42 AND Y = 6 else
"110111011111" when X = 43 AND Y = 6 else
"110111011111" when X = 44 AND Y = 6 else
"110111011111" when X = 45 AND Y = 6 else
"110111011111" when X = 46 AND Y = 6 else
"110111011111" when X = 47 AND Y = 6 else
"110111011111" when X = 48 AND Y = 6 else
"110111011111" when X = 49 AND Y = 6 else
"110111011111" when X = 50 AND Y = 6 else
"110111011111" when X = 51 AND Y = 6 else
"110111011111" when X = 52 AND Y = 6 else
"110111011111" when X = 53 AND Y = 6 else
"110111011111" when X = 54 AND Y = 6 else
"110111011111" when X = 55 AND Y = 6 else
"110111011111" when X = 56 AND Y = 6 else
"110111011111" when X = 57 AND Y = 6 else
"110111011111" when X = 58 AND Y = 6 else
"110111011111" when X = 59 AND Y = 6 else
"110111011111" when X = 60 AND Y = 6 else
"110111011111" when X = 61 AND Y = 6 else
"110111011111" when X = 62 AND Y = 6 else
"110111011111" when X = 63 AND Y = 6 else
"110111011111" when X = 64 AND Y = 6 else
"110111011111" when X = 65 AND Y = 6 else
"110111011111" when X = 66 AND Y = 6 else
"110111011111" when X = 67 AND Y = 6 else
"110111011111" when X = 68 AND Y = 6 else
"110111011111" when X = 69 AND Y = 6 else
"110111011111" when X = 70 AND Y = 6 else
"110111011111" when X = 71 AND Y = 6 else
"110111011111" when X = 72 AND Y = 6 else
"110111011111" when X = 73 AND Y = 6 else
"110111011111" when X = 74 AND Y = 6 else
"111111111111" when X = 75 AND Y = 6 else
"111111111111" when X = 76 AND Y = 6 else
"111111111111" when X = 77 AND Y = 6 else
"111111111111" when X = 78 AND Y = 6 else
"111111111111" when X = 79 AND Y = 6 else
"111111111111" when X = 80 AND Y = 6 else
"111111111111" when X = 81 AND Y = 6 else
"111111111111" when X = 82 AND Y = 6 else
"111111111111" when X = 83 AND Y = 6 else
"111111111111" when X = 84 AND Y = 6 else
"111111111111" when X = 85 AND Y = 6 else
"111111111111" when X = 86 AND Y = 6 else
"111111111111" when X = 87 AND Y = 6 else
"111111111111" when X = 88 AND Y = 6 else
"111111111111" when X = 89 AND Y = 6 else
"111111111111" when X = 90 AND Y = 6 else
"111111111111" when X = 91 AND Y = 6 else
"111111111111" when X = 92 AND Y = 6 else
"111111111111" when X = 93 AND Y = 6 else
"111111111111" when X = 94 AND Y = 6 else
"111111111111" when X = 95 AND Y = 6 else
"111111111111" when X = 96 AND Y = 6 else
"111111111111" when X = 97 AND Y = 6 else
"111111111111" when X = 98 AND Y = 6 else
"111111111111" when X = 99 AND Y = 6 else
"111111111111" when X = 100 AND Y = 6 else
"111111111111" when X = 101 AND Y = 6 else
"111111111111" when X = 102 AND Y = 6 else
"111111111111" when X = 103 AND Y = 6 else
"111111111111" when X = 104 AND Y = 6 else
"111111111111" when X = 105 AND Y = 6 else
"111111111111" when X = 106 AND Y = 6 else
"111111111111" when X = 107 AND Y = 6 else
"111111111111" when X = 108 AND Y = 6 else
"111111111111" when X = 109 AND Y = 6 else
"111111111111" when X = 110 AND Y = 6 else
"111111111111" when X = 111 AND Y = 6 else
"111111111111" when X = 112 AND Y = 6 else
"111111111111" when X = 113 AND Y = 6 else
"111111111111" when X = 114 AND Y = 6 else
"111111111111" when X = 115 AND Y = 6 else
"111111111111" when X = 116 AND Y = 6 else
"111111111111" when X = 117 AND Y = 6 else
"111111111111" when X = 118 AND Y = 6 else
"111111111111" when X = 119 AND Y = 6 else
"111111111111" when X = 120 AND Y = 6 else
"111111111111" when X = 121 AND Y = 6 else
"111111111111" when X = 122 AND Y = 6 else
"111111111111" when X = 123 AND Y = 6 else
"111111111111" when X = 124 AND Y = 6 else
"111111111111" when X = 125 AND Y = 6 else
"111111111111" when X = 126 AND Y = 6 else
"111111111111" when X = 127 AND Y = 6 else
"111111111111" when X = 128 AND Y = 6 else
"111111111111" when X = 129 AND Y = 6 else
"111111111111" when X = 130 AND Y = 6 else
"111111111111" when X = 131 AND Y = 6 else
"111111111111" when X = 132 AND Y = 6 else
"111111111111" when X = 133 AND Y = 6 else
"111111111111" when X = 134 AND Y = 6 else
"111111111111" when X = 135 AND Y = 6 else
"111111111111" when X = 136 AND Y = 6 else
"111111111111" when X = 137 AND Y = 6 else
"111111111111" when X = 138 AND Y = 6 else
"111111111111" when X = 139 AND Y = 6 else
"111111111111" when X = 140 AND Y = 6 else
"111111111111" when X = 141 AND Y = 6 else
"111111111111" when X = 142 AND Y = 6 else
"111111111111" when X = 143 AND Y = 6 else
"111111111111" when X = 144 AND Y = 6 else
"000000000000" when X = 145 AND Y = 6 else
"000000000000" when X = 146 AND Y = 6 else
"000000000000" when X = 147 AND Y = 6 else
"000000000000" when X = 148 AND Y = 6 else
"000000000000" when X = 149 AND Y = 6 else
"000000000000" when X = 150 AND Y = 6 else
"000000000000" when X = 151 AND Y = 6 else
"000000000000" when X = 152 AND Y = 6 else
"000000000000" when X = 153 AND Y = 6 else
"000000000000" when X = 154 AND Y = 6 else
"000000000000" when X = 155 AND Y = 6 else
"000000000000" when X = 156 AND Y = 6 else
"000000000000" when X = 157 AND Y = 6 else
"000000000000" when X = 158 AND Y = 6 else
"000000000000" when X = 159 AND Y = 6 else
"000000000000" when X = 160 AND Y = 6 else
"000000000000" when X = 161 AND Y = 6 else
"000000000000" when X = 162 AND Y = 6 else
"000000000000" when X = 163 AND Y = 6 else
"000000000000" when X = 164 AND Y = 6 else
"000000000000" when X = 165 AND Y = 6 else
"000000000000" when X = 166 AND Y = 6 else
"000000000000" when X = 167 AND Y = 6 else
"000000000000" when X = 168 AND Y = 6 else
"000000000000" when X = 169 AND Y = 6 else
"000000000000" when X = 170 AND Y = 6 else
"000000000000" when X = 171 AND Y = 6 else
"000000000000" when X = 172 AND Y = 6 else
"000000000000" when X = 173 AND Y = 6 else
"000000000000" when X = 174 AND Y = 6 else
"000000000000" when X = 175 AND Y = 6 else
"000000000000" when X = 176 AND Y = 6 else
"000000000000" when X = 177 AND Y = 6 else
"000000000000" when X = 178 AND Y = 6 else
"000000000000" when X = 179 AND Y = 6 else
"000000000000" when X = 180 AND Y = 6 else
"000000000000" when X = 181 AND Y = 6 else
"000000000000" when X = 182 AND Y = 6 else
"000000000000" when X = 183 AND Y = 6 else
"000000000000" when X = 184 AND Y = 6 else
"000000000000" when X = 185 AND Y = 6 else
"000000000000" when X = 186 AND Y = 6 else
"000000000000" when X = 187 AND Y = 6 else
"000000000000" when X = 188 AND Y = 6 else
"000000000000" when X = 189 AND Y = 6 else
"000000000000" when X = 190 AND Y = 6 else
"000000000000" when X = 191 AND Y = 6 else
"000000000000" when X = 192 AND Y = 6 else
"000000000000" when X = 193 AND Y = 6 else
"000000000000" when X = 194 AND Y = 6 else
"000000000000" when X = 195 AND Y = 6 else
"000000000000" when X = 196 AND Y = 6 else
"000000000000" when X = 197 AND Y = 6 else
"000000000000" when X = 198 AND Y = 6 else
"000000000000" when X = 199 AND Y = 6 else
"000000000000" when X = 200 AND Y = 6 else
"000000000000" when X = 201 AND Y = 6 else
"000000000000" when X = 202 AND Y = 6 else
"000000000000" when X = 203 AND Y = 6 else
"000000000000" when X = 204 AND Y = 6 else
"000000000000" when X = 205 AND Y = 6 else
"000000000000" when X = 206 AND Y = 6 else
"000000000000" when X = 207 AND Y = 6 else
"000000000000" when X = 208 AND Y = 6 else
"000000000000" when X = 209 AND Y = 6 else
"000000000000" when X = 210 AND Y = 6 else
"000000000000" when X = 211 AND Y = 6 else
"000000000000" when X = 212 AND Y = 6 else
"000000000000" when X = 213 AND Y = 6 else
"000000000000" when X = 214 AND Y = 6 else
"000000000000" when X = 215 AND Y = 6 else
"000000000000" when X = 216 AND Y = 6 else
"000000000000" when X = 217 AND Y = 6 else
"000000000000" when X = 218 AND Y = 6 else
"000000000000" when X = 219 AND Y = 6 else
"000000000000" when X = 220 AND Y = 6 else
"000000000000" when X = 221 AND Y = 6 else
"000000000000" when X = 222 AND Y = 6 else
"000000000000" when X = 223 AND Y = 6 else
"000000000000" when X = 224 AND Y = 6 else
"000000000000" when X = 225 AND Y = 6 else
"000000000000" when X = 226 AND Y = 6 else
"000000000000" when X = 227 AND Y = 6 else
"000000000000" when X = 228 AND Y = 6 else
"000000000000" when X = 229 AND Y = 6 else
"000000000000" when X = 230 AND Y = 6 else
"000000000000" when X = 231 AND Y = 6 else
"000000000000" when X = 232 AND Y = 6 else
"000000000000" when X = 233 AND Y = 6 else
"000000000000" when X = 234 AND Y = 6 else
"000000000000" when X = 235 AND Y = 6 else
"000000000000" when X = 236 AND Y = 6 else
"000000000000" when X = 237 AND Y = 6 else
"000000000000" when X = 238 AND Y = 6 else
"000000000000" when X = 239 AND Y = 6 else
"000000000000" when X = 240 AND Y = 6 else
"000000000000" when X = 241 AND Y = 6 else
"000000000000" when X = 242 AND Y = 6 else
"000000000000" when X = 243 AND Y = 6 else
"000000000000" when X = 244 AND Y = 6 else
"000000000000" when X = 245 AND Y = 6 else
"000000000000" when X = 246 AND Y = 6 else
"000000000000" when X = 247 AND Y = 6 else
"000000000000" when X = 248 AND Y = 6 else
"000000000000" when X = 249 AND Y = 6 else
"000000000000" when X = 250 AND Y = 6 else
"000000000000" when X = 251 AND Y = 6 else
"000000000000" when X = 252 AND Y = 6 else
"000000000000" when X = 253 AND Y = 6 else
"000000000000" when X = 254 AND Y = 6 else
"000000000000" when X = 255 AND Y = 6 else
"000000000000" when X = 256 AND Y = 6 else
"000000000000" when X = 257 AND Y = 6 else
"000000000000" when X = 258 AND Y = 6 else
"000000000000" when X = 259 AND Y = 6 else
"000000000000" when X = 260 AND Y = 6 else
"000000000000" when X = 261 AND Y = 6 else
"000000000000" when X = 262 AND Y = 6 else
"000000000000" when X = 263 AND Y = 6 else
"000000000000" when X = 264 AND Y = 6 else
"000000000000" when X = 265 AND Y = 6 else
"000000000000" when X = 266 AND Y = 6 else
"000000000000" when X = 267 AND Y = 6 else
"000000000000" when X = 268 AND Y = 6 else
"000000000000" when X = 269 AND Y = 6 else
"000000000000" when X = 270 AND Y = 6 else
"000000000000" when X = 271 AND Y = 6 else
"000000000000" when X = 272 AND Y = 6 else
"000000000000" when X = 273 AND Y = 6 else
"000000000000" when X = 274 AND Y = 6 else
"000000000000" when X = 275 AND Y = 6 else
"000000000000" when X = 276 AND Y = 6 else
"000000000000" when X = 277 AND Y = 6 else
"000000000000" when X = 278 AND Y = 6 else
"000000000000" when X = 279 AND Y = 6 else
"000000000000" when X = 280 AND Y = 6 else
"000000000000" when X = 281 AND Y = 6 else
"000000000000" when X = 282 AND Y = 6 else
"000000000000" when X = 283 AND Y = 6 else
"000000000000" when X = 284 AND Y = 6 else
"000000000000" when X = 285 AND Y = 6 else
"000000000000" when X = 286 AND Y = 6 else
"000000000000" when X = 287 AND Y = 6 else
"000000000000" when X = 288 AND Y = 6 else
"000000000000" when X = 289 AND Y = 6 else
"000000000000" when X = 290 AND Y = 6 else
"000000000000" when X = 291 AND Y = 6 else
"000000000000" when X = 292 AND Y = 6 else
"000000000000" when X = 293 AND Y = 6 else
"000000000000" when X = 294 AND Y = 6 else
"000000000000" when X = 295 AND Y = 6 else
"000000000000" when X = 296 AND Y = 6 else
"000000000000" when X = 297 AND Y = 6 else
"000000000000" when X = 298 AND Y = 6 else
"000000000000" when X = 299 AND Y = 6 else
"000000000000" when X = 300 AND Y = 6 else
"000000000000" when X = 301 AND Y = 6 else
"000000000000" when X = 302 AND Y = 6 else
"000000000000" when X = 303 AND Y = 6 else
"000000000000" when X = 304 AND Y = 6 else
"000000000000" when X = 305 AND Y = 6 else
"000000000000" when X = 306 AND Y = 6 else
"000000000000" when X = 307 AND Y = 6 else
"000000000000" when X = 308 AND Y = 6 else
"000000000000" when X = 309 AND Y = 6 else
"000000000000" when X = 310 AND Y = 6 else
"000000000000" when X = 311 AND Y = 6 else
"000000000000" when X = 312 AND Y = 6 else
"000000000000" when X = 313 AND Y = 6 else
"000000000000" when X = 314 AND Y = 6 else
"000000000000" when X = 315 AND Y = 6 else
"000000000000" when X = 316 AND Y = 6 else
"000000000000" when X = 317 AND Y = 6 else
"000000000000" when X = 318 AND Y = 6 else
"000000000000" when X = 319 AND Y = 6 else
"000000000000" when X = 320 AND Y = 6 else
"000000000000" when X = 321 AND Y = 6 else
"000000000000" when X = 322 AND Y = 6 else
"000000000000" when X = 323 AND Y = 6 else
"000000000000" when X = 324 AND Y = 6 else
"000000000000" when X = 0 AND Y = 7 else
"000000000000" when X = 1 AND Y = 7 else
"000000000000" when X = 2 AND Y = 7 else
"000000000000" when X = 3 AND Y = 7 else
"000000000000" when X = 4 AND Y = 7 else
"000000000000" when X = 5 AND Y = 7 else
"000000000000" when X = 6 AND Y = 7 else
"000000000000" when X = 7 AND Y = 7 else
"000000000000" when X = 8 AND Y = 7 else
"000000000000" when X = 9 AND Y = 7 else
"000000000000" when X = 10 AND Y = 7 else
"000000000000" when X = 11 AND Y = 7 else
"000000000000" when X = 12 AND Y = 7 else
"000000000000" when X = 13 AND Y = 7 else
"000000000000" when X = 14 AND Y = 7 else
"000000000000" when X = 15 AND Y = 7 else
"000000000000" when X = 16 AND Y = 7 else
"000000000000" when X = 17 AND Y = 7 else
"000000000000" when X = 18 AND Y = 7 else
"000000000000" when X = 19 AND Y = 7 else
"000000000000" when X = 20 AND Y = 7 else
"000000000000" when X = 21 AND Y = 7 else
"000000000000" when X = 22 AND Y = 7 else
"000000000000" when X = 23 AND Y = 7 else
"000000000000" when X = 24 AND Y = 7 else
"000000000000" when X = 25 AND Y = 7 else
"000000000000" when X = 26 AND Y = 7 else
"000000000000" when X = 27 AND Y = 7 else
"000000000000" when X = 28 AND Y = 7 else
"000000000000" when X = 29 AND Y = 7 else
"000000000000" when X = 30 AND Y = 7 else
"000000000000" when X = 31 AND Y = 7 else
"000000000000" when X = 32 AND Y = 7 else
"000000000000" when X = 33 AND Y = 7 else
"000000000000" when X = 34 AND Y = 7 else
"000000000000" when X = 35 AND Y = 7 else
"000000000000" when X = 36 AND Y = 7 else
"000000000000" when X = 37 AND Y = 7 else
"000000000000" when X = 38 AND Y = 7 else
"000000000000" when X = 39 AND Y = 7 else
"110111011111" when X = 40 AND Y = 7 else
"110111011111" when X = 41 AND Y = 7 else
"110111011111" when X = 42 AND Y = 7 else
"110111011111" when X = 43 AND Y = 7 else
"110111011111" when X = 44 AND Y = 7 else
"110111011111" when X = 45 AND Y = 7 else
"110111011111" when X = 46 AND Y = 7 else
"110111011111" when X = 47 AND Y = 7 else
"110111011111" when X = 48 AND Y = 7 else
"110111011111" when X = 49 AND Y = 7 else
"110111011111" when X = 50 AND Y = 7 else
"110111011111" when X = 51 AND Y = 7 else
"110111011111" when X = 52 AND Y = 7 else
"110111011111" when X = 53 AND Y = 7 else
"110111011111" when X = 54 AND Y = 7 else
"110111011111" when X = 55 AND Y = 7 else
"110111011111" when X = 56 AND Y = 7 else
"110111011111" when X = 57 AND Y = 7 else
"110111011111" when X = 58 AND Y = 7 else
"110111011111" when X = 59 AND Y = 7 else
"110111011111" when X = 60 AND Y = 7 else
"110111011111" when X = 61 AND Y = 7 else
"110111011111" when X = 62 AND Y = 7 else
"110111011111" when X = 63 AND Y = 7 else
"110111011111" when X = 64 AND Y = 7 else
"110111011111" when X = 65 AND Y = 7 else
"110111011111" when X = 66 AND Y = 7 else
"110111011111" when X = 67 AND Y = 7 else
"110111011111" when X = 68 AND Y = 7 else
"110111011111" when X = 69 AND Y = 7 else
"110111011111" when X = 70 AND Y = 7 else
"110111011111" when X = 71 AND Y = 7 else
"110111011111" when X = 72 AND Y = 7 else
"110111011111" when X = 73 AND Y = 7 else
"110111011111" when X = 74 AND Y = 7 else
"111111111111" when X = 75 AND Y = 7 else
"111111111111" when X = 76 AND Y = 7 else
"111111111111" when X = 77 AND Y = 7 else
"111111111111" when X = 78 AND Y = 7 else
"111111111111" when X = 79 AND Y = 7 else
"111111111111" when X = 80 AND Y = 7 else
"111111111111" when X = 81 AND Y = 7 else
"111111111111" when X = 82 AND Y = 7 else
"111111111111" when X = 83 AND Y = 7 else
"111111111111" when X = 84 AND Y = 7 else
"111111111111" when X = 85 AND Y = 7 else
"111111111111" when X = 86 AND Y = 7 else
"111111111111" when X = 87 AND Y = 7 else
"111111111111" when X = 88 AND Y = 7 else
"111111111111" when X = 89 AND Y = 7 else
"111111111111" when X = 90 AND Y = 7 else
"111111111111" when X = 91 AND Y = 7 else
"111111111111" when X = 92 AND Y = 7 else
"111111111111" when X = 93 AND Y = 7 else
"111111111111" when X = 94 AND Y = 7 else
"111111111111" when X = 95 AND Y = 7 else
"111111111111" when X = 96 AND Y = 7 else
"111111111111" when X = 97 AND Y = 7 else
"111111111111" when X = 98 AND Y = 7 else
"111111111111" when X = 99 AND Y = 7 else
"111111111111" when X = 100 AND Y = 7 else
"111111111111" when X = 101 AND Y = 7 else
"111111111111" when X = 102 AND Y = 7 else
"111111111111" when X = 103 AND Y = 7 else
"111111111111" when X = 104 AND Y = 7 else
"111111111111" when X = 105 AND Y = 7 else
"111111111111" when X = 106 AND Y = 7 else
"111111111111" when X = 107 AND Y = 7 else
"111111111111" when X = 108 AND Y = 7 else
"111111111111" when X = 109 AND Y = 7 else
"111111111111" when X = 110 AND Y = 7 else
"111111111111" when X = 111 AND Y = 7 else
"111111111111" when X = 112 AND Y = 7 else
"111111111111" when X = 113 AND Y = 7 else
"111111111111" when X = 114 AND Y = 7 else
"111111111111" when X = 115 AND Y = 7 else
"111111111111" when X = 116 AND Y = 7 else
"111111111111" when X = 117 AND Y = 7 else
"111111111111" when X = 118 AND Y = 7 else
"111111111111" when X = 119 AND Y = 7 else
"111111111111" when X = 120 AND Y = 7 else
"111111111111" when X = 121 AND Y = 7 else
"111111111111" when X = 122 AND Y = 7 else
"111111111111" when X = 123 AND Y = 7 else
"111111111111" when X = 124 AND Y = 7 else
"111111111111" when X = 125 AND Y = 7 else
"111111111111" when X = 126 AND Y = 7 else
"111111111111" when X = 127 AND Y = 7 else
"111111111111" when X = 128 AND Y = 7 else
"111111111111" when X = 129 AND Y = 7 else
"111111111111" when X = 130 AND Y = 7 else
"111111111111" when X = 131 AND Y = 7 else
"111111111111" when X = 132 AND Y = 7 else
"111111111111" when X = 133 AND Y = 7 else
"111111111111" when X = 134 AND Y = 7 else
"111111111111" when X = 135 AND Y = 7 else
"111111111111" when X = 136 AND Y = 7 else
"111111111111" when X = 137 AND Y = 7 else
"111111111111" when X = 138 AND Y = 7 else
"111111111111" when X = 139 AND Y = 7 else
"111111111111" when X = 140 AND Y = 7 else
"111111111111" when X = 141 AND Y = 7 else
"111111111111" when X = 142 AND Y = 7 else
"111111111111" when X = 143 AND Y = 7 else
"111111111111" when X = 144 AND Y = 7 else
"000000000000" when X = 145 AND Y = 7 else
"000000000000" when X = 146 AND Y = 7 else
"000000000000" when X = 147 AND Y = 7 else
"000000000000" when X = 148 AND Y = 7 else
"000000000000" when X = 149 AND Y = 7 else
"000000000000" when X = 150 AND Y = 7 else
"000000000000" when X = 151 AND Y = 7 else
"000000000000" when X = 152 AND Y = 7 else
"000000000000" when X = 153 AND Y = 7 else
"000000000000" when X = 154 AND Y = 7 else
"000000000000" when X = 155 AND Y = 7 else
"000000000000" when X = 156 AND Y = 7 else
"000000000000" when X = 157 AND Y = 7 else
"000000000000" when X = 158 AND Y = 7 else
"000000000000" when X = 159 AND Y = 7 else
"000000000000" when X = 160 AND Y = 7 else
"000000000000" when X = 161 AND Y = 7 else
"000000000000" when X = 162 AND Y = 7 else
"000000000000" when X = 163 AND Y = 7 else
"000000000000" when X = 164 AND Y = 7 else
"000000000000" when X = 165 AND Y = 7 else
"000000000000" when X = 166 AND Y = 7 else
"000000000000" when X = 167 AND Y = 7 else
"000000000000" when X = 168 AND Y = 7 else
"000000000000" when X = 169 AND Y = 7 else
"000000000000" when X = 170 AND Y = 7 else
"000000000000" when X = 171 AND Y = 7 else
"000000000000" when X = 172 AND Y = 7 else
"000000000000" when X = 173 AND Y = 7 else
"000000000000" when X = 174 AND Y = 7 else
"000000000000" when X = 175 AND Y = 7 else
"000000000000" when X = 176 AND Y = 7 else
"000000000000" when X = 177 AND Y = 7 else
"000000000000" when X = 178 AND Y = 7 else
"000000000000" when X = 179 AND Y = 7 else
"000000000000" when X = 180 AND Y = 7 else
"000000000000" when X = 181 AND Y = 7 else
"000000000000" when X = 182 AND Y = 7 else
"000000000000" when X = 183 AND Y = 7 else
"000000000000" when X = 184 AND Y = 7 else
"000000000000" when X = 185 AND Y = 7 else
"000000000000" when X = 186 AND Y = 7 else
"000000000000" when X = 187 AND Y = 7 else
"000000000000" when X = 188 AND Y = 7 else
"000000000000" when X = 189 AND Y = 7 else
"000000000000" when X = 190 AND Y = 7 else
"000000000000" when X = 191 AND Y = 7 else
"000000000000" when X = 192 AND Y = 7 else
"000000000000" when X = 193 AND Y = 7 else
"000000000000" when X = 194 AND Y = 7 else
"000000000000" when X = 195 AND Y = 7 else
"000000000000" when X = 196 AND Y = 7 else
"000000000000" when X = 197 AND Y = 7 else
"000000000000" when X = 198 AND Y = 7 else
"000000000000" when X = 199 AND Y = 7 else
"000000000000" when X = 200 AND Y = 7 else
"000000000000" when X = 201 AND Y = 7 else
"000000000000" when X = 202 AND Y = 7 else
"000000000000" when X = 203 AND Y = 7 else
"000000000000" when X = 204 AND Y = 7 else
"000000000000" when X = 205 AND Y = 7 else
"000000000000" when X = 206 AND Y = 7 else
"000000000000" when X = 207 AND Y = 7 else
"000000000000" when X = 208 AND Y = 7 else
"000000000000" when X = 209 AND Y = 7 else
"000000000000" when X = 210 AND Y = 7 else
"000000000000" when X = 211 AND Y = 7 else
"000000000000" when X = 212 AND Y = 7 else
"000000000000" when X = 213 AND Y = 7 else
"000000000000" when X = 214 AND Y = 7 else
"000000000000" when X = 215 AND Y = 7 else
"000000000000" when X = 216 AND Y = 7 else
"000000000000" when X = 217 AND Y = 7 else
"000000000000" when X = 218 AND Y = 7 else
"000000000000" when X = 219 AND Y = 7 else
"000000000000" when X = 220 AND Y = 7 else
"000000000000" when X = 221 AND Y = 7 else
"000000000000" when X = 222 AND Y = 7 else
"000000000000" when X = 223 AND Y = 7 else
"000000000000" when X = 224 AND Y = 7 else
"000000000000" when X = 225 AND Y = 7 else
"000000000000" when X = 226 AND Y = 7 else
"000000000000" when X = 227 AND Y = 7 else
"000000000000" when X = 228 AND Y = 7 else
"000000000000" when X = 229 AND Y = 7 else
"000000000000" when X = 230 AND Y = 7 else
"000000000000" when X = 231 AND Y = 7 else
"000000000000" when X = 232 AND Y = 7 else
"000000000000" when X = 233 AND Y = 7 else
"000000000000" when X = 234 AND Y = 7 else
"000000000000" when X = 235 AND Y = 7 else
"000000000000" when X = 236 AND Y = 7 else
"000000000000" when X = 237 AND Y = 7 else
"000000000000" when X = 238 AND Y = 7 else
"000000000000" when X = 239 AND Y = 7 else
"000000000000" when X = 240 AND Y = 7 else
"000000000000" when X = 241 AND Y = 7 else
"000000000000" when X = 242 AND Y = 7 else
"000000000000" when X = 243 AND Y = 7 else
"000000000000" when X = 244 AND Y = 7 else
"000000000000" when X = 245 AND Y = 7 else
"000000000000" when X = 246 AND Y = 7 else
"000000000000" when X = 247 AND Y = 7 else
"000000000000" when X = 248 AND Y = 7 else
"000000000000" when X = 249 AND Y = 7 else
"000000000000" when X = 250 AND Y = 7 else
"000000000000" when X = 251 AND Y = 7 else
"000000000000" when X = 252 AND Y = 7 else
"000000000000" when X = 253 AND Y = 7 else
"000000000000" when X = 254 AND Y = 7 else
"000000000000" when X = 255 AND Y = 7 else
"000000000000" when X = 256 AND Y = 7 else
"000000000000" when X = 257 AND Y = 7 else
"000000000000" when X = 258 AND Y = 7 else
"000000000000" when X = 259 AND Y = 7 else
"000000000000" when X = 260 AND Y = 7 else
"000000000000" when X = 261 AND Y = 7 else
"000000000000" when X = 262 AND Y = 7 else
"000000000000" when X = 263 AND Y = 7 else
"000000000000" when X = 264 AND Y = 7 else
"000000000000" when X = 265 AND Y = 7 else
"000000000000" when X = 266 AND Y = 7 else
"000000000000" when X = 267 AND Y = 7 else
"000000000000" when X = 268 AND Y = 7 else
"000000000000" when X = 269 AND Y = 7 else
"000000000000" when X = 270 AND Y = 7 else
"000000000000" when X = 271 AND Y = 7 else
"000000000000" when X = 272 AND Y = 7 else
"000000000000" when X = 273 AND Y = 7 else
"000000000000" when X = 274 AND Y = 7 else
"000000000000" when X = 275 AND Y = 7 else
"000000000000" when X = 276 AND Y = 7 else
"000000000000" when X = 277 AND Y = 7 else
"000000000000" when X = 278 AND Y = 7 else
"000000000000" when X = 279 AND Y = 7 else
"000000000000" when X = 280 AND Y = 7 else
"000000000000" when X = 281 AND Y = 7 else
"000000000000" when X = 282 AND Y = 7 else
"000000000000" when X = 283 AND Y = 7 else
"000000000000" when X = 284 AND Y = 7 else
"000000000000" when X = 285 AND Y = 7 else
"000000000000" when X = 286 AND Y = 7 else
"000000000000" when X = 287 AND Y = 7 else
"000000000000" when X = 288 AND Y = 7 else
"000000000000" when X = 289 AND Y = 7 else
"000000000000" when X = 290 AND Y = 7 else
"000000000000" when X = 291 AND Y = 7 else
"000000000000" when X = 292 AND Y = 7 else
"000000000000" when X = 293 AND Y = 7 else
"000000000000" when X = 294 AND Y = 7 else
"000000000000" when X = 295 AND Y = 7 else
"000000000000" when X = 296 AND Y = 7 else
"000000000000" when X = 297 AND Y = 7 else
"000000000000" when X = 298 AND Y = 7 else
"000000000000" when X = 299 AND Y = 7 else
"000000000000" when X = 300 AND Y = 7 else
"000000000000" when X = 301 AND Y = 7 else
"000000000000" when X = 302 AND Y = 7 else
"000000000000" when X = 303 AND Y = 7 else
"000000000000" when X = 304 AND Y = 7 else
"000000000000" when X = 305 AND Y = 7 else
"000000000000" when X = 306 AND Y = 7 else
"000000000000" when X = 307 AND Y = 7 else
"000000000000" when X = 308 AND Y = 7 else
"000000000000" when X = 309 AND Y = 7 else
"000000000000" when X = 310 AND Y = 7 else
"000000000000" when X = 311 AND Y = 7 else
"000000000000" when X = 312 AND Y = 7 else
"000000000000" when X = 313 AND Y = 7 else
"000000000000" when X = 314 AND Y = 7 else
"000000000000" when X = 315 AND Y = 7 else
"000000000000" when X = 316 AND Y = 7 else
"000000000000" when X = 317 AND Y = 7 else
"000000000000" when X = 318 AND Y = 7 else
"000000000000" when X = 319 AND Y = 7 else
"000000000000" when X = 320 AND Y = 7 else
"000000000000" when X = 321 AND Y = 7 else
"000000000000" when X = 322 AND Y = 7 else
"000000000000" when X = 323 AND Y = 7 else
"000000000000" when X = 324 AND Y = 7 else
"000000000000" when X = 0 AND Y = 8 else
"000000000000" when X = 1 AND Y = 8 else
"000000000000" when X = 2 AND Y = 8 else
"000000000000" when X = 3 AND Y = 8 else
"000000000000" when X = 4 AND Y = 8 else
"000000000000" when X = 5 AND Y = 8 else
"000000000000" when X = 6 AND Y = 8 else
"000000000000" when X = 7 AND Y = 8 else
"000000000000" when X = 8 AND Y = 8 else
"000000000000" when X = 9 AND Y = 8 else
"000000000000" when X = 10 AND Y = 8 else
"000000000000" when X = 11 AND Y = 8 else
"000000000000" when X = 12 AND Y = 8 else
"000000000000" when X = 13 AND Y = 8 else
"000000000000" when X = 14 AND Y = 8 else
"000000000000" when X = 15 AND Y = 8 else
"000000000000" when X = 16 AND Y = 8 else
"000000000000" when X = 17 AND Y = 8 else
"000000000000" when X = 18 AND Y = 8 else
"000000000000" when X = 19 AND Y = 8 else
"000000000000" when X = 20 AND Y = 8 else
"000000000000" when X = 21 AND Y = 8 else
"000000000000" when X = 22 AND Y = 8 else
"000000000000" when X = 23 AND Y = 8 else
"000000000000" when X = 24 AND Y = 8 else
"000000000000" when X = 25 AND Y = 8 else
"000000000000" when X = 26 AND Y = 8 else
"000000000000" when X = 27 AND Y = 8 else
"000000000000" when X = 28 AND Y = 8 else
"000000000000" when X = 29 AND Y = 8 else
"000000000000" when X = 30 AND Y = 8 else
"000000000000" when X = 31 AND Y = 8 else
"000000000000" when X = 32 AND Y = 8 else
"000000000000" when X = 33 AND Y = 8 else
"000000000000" when X = 34 AND Y = 8 else
"000000000000" when X = 35 AND Y = 8 else
"000000000000" when X = 36 AND Y = 8 else
"000000000000" when X = 37 AND Y = 8 else
"000000000000" when X = 38 AND Y = 8 else
"000000000000" when X = 39 AND Y = 8 else
"110111011111" when X = 40 AND Y = 8 else
"110111011111" when X = 41 AND Y = 8 else
"110111011111" when X = 42 AND Y = 8 else
"110111011111" when X = 43 AND Y = 8 else
"110111011111" when X = 44 AND Y = 8 else
"110111011111" when X = 45 AND Y = 8 else
"110111011111" when X = 46 AND Y = 8 else
"110111011111" when X = 47 AND Y = 8 else
"110111011111" when X = 48 AND Y = 8 else
"110111011111" when X = 49 AND Y = 8 else
"110111011111" when X = 50 AND Y = 8 else
"110111011111" when X = 51 AND Y = 8 else
"110111011111" when X = 52 AND Y = 8 else
"110111011111" when X = 53 AND Y = 8 else
"110111011111" when X = 54 AND Y = 8 else
"110111011111" when X = 55 AND Y = 8 else
"110111011111" when X = 56 AND Y = 8 else
"110111011111" when X = 57 AND Y = 8 else
"110111011111" when X = 58 AND Y = 8 else
"110111011111" when X = 59 AND Y = 8 else
"110111011111" when X = 60 AND Y = 8 else
"110111011111" when X = 61 AND Y = 8 else
"110111011111" when X = 62 AND Y = 8 else
"110111011111" when X = 63 AND Y = 8 else
"110111011111" when X = 64 AND Y = 8 else
"110111011111" when X = 65 AND Y = 8 else
"110111011111" when X = 66 AND Y = 8 else
"110111011111" when X = 67 AND Y = 8 else
"110111011111" when X = 68 AND Y = 8 else
"110111011111" when X = 69 AND Y = 8 else
"110111011111" when X = 70 AND Y = 8 else
"110111011111" when X = 71 AND Y = 8 else
"110111011111" when X = 72 AND Y = 8 else
"110111011111" when X = 73 AND Y = 8 else
"110111011111" when X = 74 AND Y = 8 else
"111111111111" when X = 75 AND Y = 8 else
"111111111111" when X = 76 AND Y = 8 else
"111111111111" when X = 77 AND Y = 8 else
"111111111111" when X = 78 AND Y = 8 else
"111111111111" when X = 79 AND Y = 8 else
"111111111111" when X = 80 AND Y = 8 else
"111111111111" when X = 81 AND Y = 8 else
"111111111111" when X = 82 AND Y = 8 else
"111111111111" when X = 83 AND Y = 8 else
"111111111111" when X = 84 AND Y = 8 else
"111111111111" when X = 85 AND Y = 8 else
"111111111111" when X = 86 AND Y = 8 else
"111111111111" when X = 87 AND Y = 8 else
"111111111111" when X = 88 AND Y = 8 else
"111111111111" when X = 89 AND Y = 8 else
"111111111111" when X = 90 AND Y = 8 else
"111111111111" when X = 91 AND Y = 8 else
"111111111111" when X = 92 AND Y = 8 else
"111111111111" when X = 93 AND Y = 8 else
"111111111111" when X = 94 AND Y = 8 else
"111111111111" when X = 95 AND Y = 8 else
"111111111111" when X = 96 AND Y = 8 else
"111111111111" when X = 97 AND Y = 8 else
"111111111111" when X = 98 AND Y = 8 else
"111111111111" when X = 99 AND Y = 8 else
"111111111111" when X = 100 AND Y = 8 else
"111111111111" when X = 101 AND Y = 8 else
"111111111111" when X = 102 AND Y = 8 else
"111111111111" when X = 103 AND Y = 8 else
"111111111111" when X = 104 AND Y = 8 else
"111111111111" when X = 105 AND Y = 8 else
"111111111111" when X = 106 AND Y = 8 else
"111111111111" when X = 107 AND Y = 8 else
"111111111111" when X = 108 AND Y = 8 else
"111111111111" when X = 109 AND Y = 8 else
"111111111111" when X = 110 AND Y = 8 else
"111111111111" when X = 111 AND Y = 8 else
"111111111111" when X = 112 AND Y = 8 else
"111111111111" when X = 113 AND Y = 8 else
"111111111111" when X = 114 AND Y = 8 else
"111111111111" when X = 115 AND Y = 8 else
"111111111111" when X = 116 AND Y = 8 else
"111111111111" when X = 117 AND Y = 8 else
"111111111111" when X = 118 AND Y = 8 else
"111111111111" when X = 119 AND Y = 8 else
"111111111111" when X = 120 AND Y = 8 else
"111111111111" when X = 121 AND Y = 8 else
"111111111111" when X = 122 AND Y = 8 else
"111111111111" when X = 123 AND Y = 8 else
"111111111111" when X = 124 AND Y = 8 else
"111111111111" when X = 125 AND Y = 8 else
"111111111111" when X = 126 AND Y = 8 else
"111111111111" when X = 127 AND Y = 8 else
"111111111111" when X = 128 AND Y = 8 else
"111111111111" when X = 129 AND Y = 8 else
"111111111111" when X = 130 AND Y = 8 else
"111111111111" when X = 131 AND Y = 8 else
"111111111111" when X = 132 AND Y = 8 else
"111111111111" when X = 133 AND Y = 8 else
"111111111111" when X = 134 AND Y = 8 else
"111111111111" when X = 135 AND Y = 8 else
"111111111111" when X = 136 AND Y = 8 else
"111111111111" when X = 137 AND Y = 8 else
"111111111111" when X = 138 AND Y = 8 else
"111111111111" when X = 139 AND Y = 8 else
"111111111111" when X = 140 AND Y = 8 else
"111111111111" when X = 141 AND Y = 8 else
"111111111111" when X = 142 AND Y = 8 else
"111111111111" when X = 143 AND Y = 8 else
"111111111111" when X = 144 AND Y = 8 else
"000000000000" when X = 145 AND Y = 8 else
"000000000000" when X = 146 AND Y = 8 else
"000000000000" when X = 147 AND Y = 8 else
"000000000000" when X = 148 AND Y = 8 else
"000000000000" when X = 149 AND Y = 8 else
"000000000000" when X = 150 AND Y = 8 else
"000000000000" when X = 151 AND Y = 8 else
"000000000000" when X = 152 AND Y = 8 else
"000000000000" when X = 153 AND Y = 8 else
"000000000000" when X = 154 AND Y = 8 else
"000000000000" when X = 155 AND Y = 8 else
"000000000000" when X = 156 AND Y = 8 else
"000000000000" when X = 157 AND Y = 8 else
"000000000000" when X = 158 AND Y = 8 else
"000000000000" when X = 159 AND Y = 8 else
"000000000000" when X = 160 AND Y = 8 else
"000000000000" when X = 161 AND Y = 8 else
"000000000000" when X = 162 AND Y = 8 else
"000000000000" when X = 163 AND Y = 8 else
"000000000000" when X = 164 AND Y = 8 else
"000000000000" when X = 165 AND Y = 8 else
"000000000000" when X = 166 AND Y = 8 else
"000000000000" when X = 167 AND Y = 8 else
"000000000000" when X = 168 AND Y = 8 else
"000000000000" when X = 169 AND Y = 8 else
"000000000000" when X = 170 AND Y = 8 else
"000000000000" when X = 171 AND Y = 8 else
"000000000000" when X = 172 AND Y = 8 else
"000000000000" when X = 173 AND Y = 8 else
"000000000000" when X = 174 AND Y = 8 else
"000000000000" when X = 175 AND Y = 8 else
"000000000000" when X = 176 AND Y = 8 else
"000000000000" when X = 177 AND Y = 8 else
"000000000000" when X = 178 AND Y = 8 else
"000000000000" when X = 179 AND Y = 8 else
"000000000000" when X = 180 AND Y = 8 else
"000000000000" when X = 181 AND Y = 8 else
"000000000000" when X = 182 AND Y = 8 else
"000000000000" when X = 183 AND Y = 8 else
"000000000000" when X = 184 AND Y = 8 else
"000000000000" when X = 185 AND Y = 8 else
"000000000000" when X = 186 AND Y = 8 else
"000000000000" when X = 187 AND Y = 8 else
"000000000000" when X = 188 AND Y = 8 else
"000000000000" when X = 189 AND Y = 8 else
"000000000000" when X = 190 AND Y = 8 else
"000000000000" when X = 191 AND Y = 8 else
"000000000000" when X = 192 AND Y = 8 else
"000000000000" when X = 193 AND Y = 8 else
"000000000000" when X = 194 AND Y = 8 else
"000000000000" when X = 195 AND Y = 8 else
"000000000000" when X = 196 AND Y = 8 else
"000000000000" when X = 197 AND Y = 8 else
"000000000000" when X = 198 AND Y = 8 else
"000000000000" when X = 199 AND Y = 8 else
"000000000000" when X = 200 AND Y = 8 else
"000000000000" when X = 201 AND Y = 8 else
"000000000000" when X = 202 AND Y = 8 else
"000000000000" when X = 203 AND Y = 8 else
"000000000000" when X = 204 AND Y = 8 else
"000000000000" when X = 205 AND Y = 8 else
"000000000000" when X = 206 AND Y = 8 else
"000000000000" when X = 207 AND Y = 8 else
"000000000000" when X = 208 AND Y = 8 else
"000000000000" when X = 209 AND Y = 8 else
"000000000000" when X = 210 AND Y = 8 else
"000000000000" when X = 211 AND Y = 8 else
"000000000000" when X = 212 AND Y = 8 else
"000000000000" when X = 213 AND Y = 8 else
"000000000000" when X = 214 AND Y = 8 else
"000000000000" when X = 215 AND Y = 8 else
"000000000000" when X = 216 AND Y = 8 else
"000000000000" when X = 217 AND Y = 8 else
"000000000000" when X = 218 AND Y = 8 else
"000000000000" when X = 219 AND Y = 8 else
"000000000000" when X = 220 AND Y = 8 else
"000000000000" when X = 221 AND Y = 8 else
"000000000000" when X = 222 AND Y = 8 else
"000000000000" when X = 223 AND Y = 8 else
"000000000000" when X = 224 AND Y = 8 else
"000000000000" when X = 225 AND Y = 8 else
"000000000000" when X = 226 AND Y = 8 else
"000000000000" when X = 227 AND Y = 8 else
"000000000000" when X = 228 AND Y = 8 else
"000000000000" when X = 229 AND Y = 8 else
"000000000000" when X = 230 AND Y = 8 else
"000000000000" when X = 231 AND Y = 8 else
"000000000000" when X = 232 AND Y = 8 else
"000000000000" when X = 233 AND Y = 8 else
"000000000000" when X = 234 AND Y = 8 else
"000000000000" when X = 235 AND Y = 8 else
"000000000000" when X = 236 AND Y = 8 else
"000000000000" when X = 237 AND Y = 8 else
"000000000000" when X = 238 AND Y = 8 else
"000000000000" when X = 239 AND Y = 8 else
"000000000000" when X = 240 AND Y = 8 else
"000000000000" when X = 241 AND Y = 8 else
"000000000000" when X = 242 AND Y = 8 else
"000000000000" when X = 243 AND Y = 8 else
"000000000000" when X = 244 AND Y = 8 else
"000000000000" when X = 245 AND Y = 8 else
"000000000000" when X = 246 AND Y = 8 else
"000000000000" when X = 247 AND Y = 8 else
"000000000000" when X = 248 AND Y = 8 else
"000000000000" when X = 249 AND Y = 8 else
"000000000000" when X = 250 AND Y = 8 else
"000000000000" when X = 251 AND Y = 8 else
"000000000000" when X = 252 AND Y = 8 else
"000000000000" when X = 253 AND Y = 8 else
"000000000000" when X = 254 AND Y = 8 else
"000000000000" when X = 255 AND Y = 8 else
"000000000000" when X = 256 AND Y = 8 else
"000000000000" when X = 257 AND Y = 8 else
"000000000000" when X = 258 AND Y = 8 else
"000000000000" when X = 259 AND Y = 8 else
"000000000000" when X = 260 AND Y = 8 else
"000000000000" when X = 261 AND Y = 8 else
"000000000000" when X = 262 AND Y = 8 else
"000000000000" when X = 263 AND Y = 8 else
"000000000000" when X = 264 AND Y = 8 else
"000000000000" when X = 265 AND Y = 8 else
"000000000000" when X = 266 AND Y = 8 else
"000000000000" when X = 267 AND Y = 8 else
"000000000000" when X = 268 AND Y = 8 else
"000000000000" when X = 269 AND Y = 8 else
"000000000000" when X = 270 AND Y = 8 else
"000000000000" when X = 271 AND Y = 8 else
"000000000000" when X = 272 AND Y = 8 else
"000000000000" when X = 273 AND Y = 8 else
"000000000000" when X = 274 AND Y = 8 else
"000000000000" when X = 275 AND Y = 8 else
"000000000000" when X = 276 AND Y = 8 else
"000000000000" when X = 277 AND Y = 8 else
"000000000000" when X = 278 AND Y = 8 else
"000000000000" when X = 279 AND Y = 8 else
"000000000000" when X = 280 AND Y = 8 else
"000000000000" when X = 281 AND Y = 8 else
"000000000000" when X = 282 AND Y = 8 else
"000000000000" when X = 283 AND Y = 8 else
"000000000000" when X = 284 AND Y = 8 else
"000000000000" when X = 285 AND Y = 8 else
"000000000000" when X = 286 AND Y = 8 else
"000000000000" when X = 287 AND Y = 8 else
"000000000000" when X = 288 AND Y = 8 else
"000000000000" when X = 289 AND Y = 8 else
"000000000000" when X = 290 AND Y = 8 else
"000000000000" when X = 291 AND Y = 8 else
"000000000000" when X = 292 AND Y = 8 else
"000000000000" when X = 293 AND Y = 8 else
"000000000000" when X = 294 AND Y = 8 else
"000000000000" when X = 295 AND Y = 8 else
"000000000000" when X = 296 AND Y = 8 else
"000000000000" when X = 297 AND Y = 8 else
"000000000000" when X = 298 AND Y = 8 else
"000000000000" when X = 299 AND Y = 8 else
"000000000000" when X = 300 AND Y = 8 else
"000000000000" when X = 301 AND Y = 8 else
"000000000000" when X = 302 AND Y = 8 else
"000000000000" when X = 303 AND Y = 8 else
"000000000000" when X = 304 AND Y = 8 else
"000000000000" when X = 305 AND Y = 8 else
"000000000000" when X = 306 AND Y = 8 else
"000000000000" when X = 307 AND Y = 8 else
"000000000000" when X = 308 AND Y = 8 else
"000000000000" when X = 309 AND Y = 8 else
"000000000000" when X = 310 AND Y = 8 else
"000000000000" when X = 311 AND Y = 8 else
"000000000000" when X = 312 AND Y = 8 else
"000000000000" when X = 313 AND Y = 8 else
"000000000000" when X = 314 AND Y = 8 else
"000000000000" when X = 315 AND Y = 8 else
"000000000000" when X = 316 AND Y = 8 else
"000000000000" when X = 317 AND Y = 8 else
"000000000000" when X = 318 AND Y = 8 else
"000000000000" when X = 319 AND Y = 8 else
"000000000000" when X = 320 AND Y = 8 else
"000000000000" when X = 321 AND Y = 8 else
"000000000000" when X = 322 AND Y = 8 else
"000000000000" when X = 323 AND Y = 8 else
"000000000000" when X = 324 AND Y = 8 else
"000000000000" when X = 0 AND Y = 9 else
"000000000000" when X = 1 AND Y = 9 else
"000000000000" when X = 2 AND Y = 9 else
"000000000000" when X = 3 AND Y = 9 else
"000000000000" when X = 4 AND Y = 9 else
"000000000000" when X = 5 AND Y = 9 else
"000000000000" when X = 6 AND Y = 9 else
"000000000000" when X = 7 AND Y = 9 else
"000000000000" when X = 8 AND Y = 9 else
"000000000000" when X = 9 AND Y = 9 else
"000000000000" when X = 10 AND Y = 9 else
"000000000000" when X = 11 AND Y = 9 else
"000000000000" when X = 12 AND Y = 9 else
"000000000000" when X = 13 AND Y = 9 else
"000000000000" when X = 14 AND Y = 9 else
"000000000000" when X = 15 AND Y = 9 else
"000000000000" when X = 16 AND Y = 9 else
"000000000000" when X = 17 AND Y = 9 else
"000000000000" when X = 18 AND Y = 9 else
"000000000000" when X = 19 AND Y = 9 else
"000000000000" when X = 20 AND Y = 9 else
"000000000000" when X = 21 AND Y = 9 else
"000000000000" when X = 22 AND Y = 9 else
"000000000000" when X = 23 AND Y = 9 else
"000000000000" when X = 24 AND Y = 9 else
"000000000000" when X = 25 AND Y = 9 else
"000000000000" when X = 26 AND Y = 9 else
"000000000000" when X = 27 AND Y = 9 else
"000000000000" when X = 28 AND Y = 9 else
"000000000000" when X = 29 AND Y = 9 else
"000000000000" when X = 30 AND Y = 9 else
"000000000000" when X = 31 AND Y = 9 else
"000000000000" when X = 32 AND Y = 9 else
"000000000000" when X = 33 AND Y = 9 else
"000000000000" when X = 34 AND Y = 9 else
"000000000000" when X = 35 AND Y = 9 else
"000000000000" when X = 36 AND Y = 9 else
"000000000000" when X = 37 AND Y = 9 else
"000000000000" when X = 38 AND Y = 9 else
"000000000000" when X = 39 AND Y = 9 else
"110111011111" when X = 40 AND Y = 9 else
"110111011111" when X = 41 AND Y = 9 else
"110111011111" when X = 42 AND Y = 9 else
"110111011111" when X = 43 AND Y = 9 else
"110111011111" when X = 44 AND Y = 9 else
"110111011111" when X = 45 AND Y = 9 else
"110111011111" when X = 46 AND Y = 9 else
"110111011111" when X = 47 AND Y = 9 else
"110111011111" when X = 48 AND Y = 9 else
"110111011111" when X = 49 AND Y = 9 else
"110111011111" when X = 50 AND Y = 9 else
"110111011111" when X = 51 AND Y = 9 else
"110111011111" when X = 52 AND Y = 9 else
"110111011111" when X = 53 AND Y = 9 else
"110111011111" when X = 54 AND Y = 9 else
"110111011111" when X = 55 AND Y = 9 else
"110111011111" when X = 56 AND Y = 9 else
"110111011111" when X = 57 AND Y = 9 else
"110111011111" when X = 58 AND Y = 9 else
"110111011111" when X = 59 AND Y = 9 else
"110111011111" when X = 60 AND Y = 9 else
"110111011111" when X = 61 AND Y = 9 else
"110111011111" when X = 62 AND Y = 9 else
"110111011111" when X = 63 AND Y = 9 else
"110111011111" when X = 64 AND Y = 9 else
"110111011111" when X = 65 AND Y = 9 else
"110111011111" when X = 66 AND Y = 9 else
"110111011111" when X = 67 AND Y = 9 else
"110111011111" when X = 68 AND Y = 9 else
"110111011111" when X = 69 AND Y = 9 else
"110111011111" when X = 70 AND Y = 9 else
"110111011111" when X = 71 AND Y = 9 else
"110111011111" when X = 72 AND Y = 9 else
"110111011111" when X = 73 AND Y = 9 else
"110111011111" when X = 74 AND Y = 9 else
"111111111111" when X = 75 AND Y = 9 else
"111111111111" when X = 76 AND Y = 9 else
"111111111111" when X = 77 AND Y = 9 else
"111111111111" when X = 78 AND Y = 9 else
"111111111111" when X = 79 AND Y = 9 else
"111111111111" when X = 80 AND Y = 9 else
"111111111111" when X = 81 AND Y = 9 else
"111111111111" when X = 82 AND Y = 9 else
"111111111111" when X = 83 AND Y = 9 else
"111111111111" when X = 84 AND Y = 9 else
"111111111111" when X = 85 AND Y = 9 else
"111111111111" when X = 86 AND Y = 9 else
"111111111111" when X = 87 AND Y = 9 else
"111111111111" when X = 88 AND Y = 9 else
"111111111111" when X = 89 AND Y = 9 else
"111111111111" when X = 90 AND Y = 9 else
"111111111111" when X = 91 AND Y = 9 else
"111111111111" when X = 92 AND Y = 9 else
"111111111111" when X = 93 AND Y = 9 else
"111111111111" when X = 94 AND Y = 9 else
"111111111111" when X = 95 AND Y = 9 else
"111111111111" when X = 96 AND Y = 9 else
"111111111111" when X = 97 AND Y = 9 else
"111111111111" when X = 98 AND Y = 9 else
"111111111111" when X = 99 AND Y = 9 else
"111111111111" when X = 100 AND Y = 9 else
"111111111111" when X = 101 AND Y = 9 else
"111111111111" when X = 102 AND Y = 9 else
"111111111111" when X = 103 AND Y = 9 else
"111111111111" when X = 104 AND Y = 9 else
"111111111111" when X = 105 AND Y = 9 else
"111111111111" when X = 106 AND Y = 9 else
"111111111111" when X = 107 AND Y = 9 else
"111111111111" when X = 108 AND Y = 9 else
"111111111111" when X = 109 AND Y = 9 else
"111111111111" when X = 110 AND Y = 9 else
"111111111111" when X = 111 AND Y = 9 else
"111111111111" when X = 112 AND Y = 9 else
"111111111111" when X = 113 AND Y = 9 else
"111111111111" when X = 114 AND Y = 9 else
"111111111111" when X = 115 AND Y = 9 else
"111111111111" when X = 116 AND Y = 9 else
"111111111111" when X = 117 AND Y = 9 else
"111111111111" when X = 118 AND Y = 9 else
"111111111111" when X = 119 AND Y = 9 else
"111111111111" when X = 120 AND Y = 9 else
"111111111111" when X = 121 AND Y = 9 else
"111111111111" when X = 122 AND Y = 9 else
"111111111111" when X = 123 AND Y = 9 else
"111111111111" when X = 124 AND Y = 9 else
"111111111111" when X = 125 AND Y = 9 else
"111111111111" when X = 126 AND Y = 9 else
"111111111111" when X = 127 AND Y = 9 else
"111111111111" when X = 128 AND Y = 9 else
"111111111111" when X = 129 AND Y = 9 else
"111111111111" when X = 130 AND Y = 9 else
"111111111111" when X = 131 AND Y = 9 else
"111111111111" when X = 132 AND Y = 9 else
"111111111111" when X = 133 AND Y = 9 else
"111111111111" when X = 134 AND Y = 9 else
"111111111111" when X = 135 AND Y = 9 else
"111111111111" when X = 136 AND Y = 9 else
"111111111111" when X = 137 AND Y = 9 else
"111111111111" when X = 138 AND Y = 9 else
"111111111111" when X = 139 AND Y = 9 else
"111111111111" when X = 140 AND Y = 9 else
"111111111111" when X = 141 AND Y = 9 else
"111111111111" when X = 142 AND Y = 9 else
"111111111111" when X = 143 AND Y = 9 else
"111111111111" when X = 144 AND Y = 9 else
"000000000000" when X = 145 AND Y = 9 else
"000000000000" when X = 146 AND Y = 9 else
"000000000000" when X = 147 AND Y = 9 else
"000000000000" when X = 148 AND Y = 9 else
"000000000000" when X = 149 AND Y = 9 else
"000000000000" when X = 150 AND Y = 9 else
"000000000000" when X = 151 AND Y = 9 else
"000000000000" when X = 152 AND Y = 9 else
"000000000000" when X = 153 AND Y = 9 else
"000000000000" when X = 154 AND Y = 9 else
"000000000000" when X = 155 AND Y = 9 else
"000000000000" when X = 156 AND Y = 9 else
"000000000000" when X = 157 AND Y = 9 else
"000000000000" when X = 158 AND Y = 9 else
"000000000000" when X = 159 AND Y = 9 else
"000000000000" when X = 160 AND Y = 9 else
"000000000000" when X = 161 AND Y = 9 else
"000000000000" when X = 162 AND Y = 9 else
"000000000000" when X = 163 AND Y = 9 else
"000000000000" when X = 164 AND Y = 9 else
"000000000000" when X = 165 AND Y = 9 else
"000000000000" when X = 166 AND Y = 9 else
"000000000000" when X = 167 AND Y = 9 else
"000000000000" when X = 168 AND Y = 9 else
"000000000000" when X = 169 AND Y = 9 else
"000000000000" when X = 170 AND Y = 9 else
"000000000000" when X = 171 AND Y = 9 else
"000000000000" when X = 172 AND Y = 9 else
"000000000000" when X = 173 AND Y = 9 else
"000000000000" when X = 174 AND Y = 9 else
"000000000000" when X = 175 AND Y = 9 else
"000000000000" when X = 176 AND Y = 9 else
"000000000000" when X = 177 AND Y = 9 else
"000000000000" when X = 178 AND Y = 9 else
"000000000000" when X = 179 AND Y = 9 else
"000000000000" when X = 180 AND Y = 9 else
"000000000000" when X = 181 AND Y = 9 else
"000000000000" when X = 182 AND Y = 9 else
"000000000000" when X = 183 AND Y = 9 else
"000000000000" when X = 184 AND Y = 9 else
"000000000000" when X = 185 AND Y = 9 else
"000000000000" when X = 186 AND Y = 9 else
"000000000000" when X = 187 AND Y = 9 else
"000000000000" when X = 188 AND Y = 9 else
"000000000000" when X = 189 AND Y = 9 else
"000000000000" when X = 190 AND Y = 9 else
"000000000000" when X = 191 AND Y = 9 else
"000000000000" when X = 192 AND Y = 9 else
"000000000000" when X = 193 AND Y = 9 else
"000000000000" when X = 194 AND Y = 9 else
"000000000000" when X = 195 AND Y = 9 else
"000000000000" when X = 196 AND Y = 9 else
"000000000000" when X = 197 AND Y = 9 else
"000000000000" when X = 198 AND Y = 9 else
"000000000000" when X = 199 AND Y = 9 else
"000000000000" when X = 200 AND Y = 9 else
"000000000000" when X = 201 AND Y = 9 else
"000000000000" when X = 202 AND Y = 9 else
"000000000000" when X = 203 AND Y = 9 else
"000000000000" when X = 204 AND Y = 9 else
"000000000000" when X = 205 AND Y = 9 else
"000000000000" when X = 206 AND Y = 9 else
"000000000000" when X = 207 AND Y = 9 else
"000000000000" when X = 208 AND Y = 9 else
"000000000000" when X = 209 AND Y = 9 else
"000000000000" when X = 210 AND Y = 9 else
"000000000000" when X = 211 AND Y = 9 else
"000000000000" when X = 212 AND Y = 9 else
"000000000000" when X = 213 AND Y = 9 else
"000000000000" when X = 214 AND Y = 9 else
"000000000000" when X = 215 AND Y = 9 else
"000000000000" when X = 216 AND Y = 9 else
"000000000000" when X = 217 AND Y = 9 else
"000000000000" when X = 218 AND Y = 9 else
"000000000000" when X = 219 AND Y = 9 else
"000000000000" when X = 220 AND Y = 9 else
"000000000000" when X = 221 AND Y = 9 else
"000000000000" when X = 222 AND Y = 9 else
"000000000000" when X = 223 AND Y = 9 else
"000000000000" when X = 224 AND Y = 9 else
"000000000000" when X = 225 AND Y = 9 else
"000000000000" when X = 226 AND Y = 9 else
"000000000000" when X = 227 AND Y = 9 else
"000000000000" when X = 228 AND Y = 9 else
"000000000000" when X = 229 AND Y = 9 else
"000000000000" when X = 230 AND Y = 9 else
"000000000000" when X = 231 AND Y = 9 else
"000000000000" when X = 232 AND Y = 9 else
"000000000000" when X = 233 AND Y = 9 else
"000000000000" when X = 234 AND Y = 9 else
"000000000000" when X = 235 AND Y = 9 else
"000000000000" when X = 236 AND Y = 9 else
"000000000000" when X = 237 AND Y = 9 else
"000000000000" when X = 238 AND Y = 9 else
"000000000000" when X = 239 AND Y = 9 else
"000000000000" when X = 240 AND Y = 9 else
"000000000000" when X = 241 AND Y = 9 else
"000000000000" when X = 242 AND Y = 9 else
"000000000000" when X = 243 AND Y = 9 else
"000000000000" when X = 244 AND Y = 9 else
"000000000000" when X = 245 AND Y = 9 else
"000000000000" when X = 246 AND Y = 9 else
"000000000000" when X = 247 AND Y = 9 else
"000000000000" when X = 248 AND Y = 9 else
"000000000000" when X = 249 AND Y = 9 else
"000000000000" when X = 250 AND Y = 9 else
"000000000000" when X = 251 AND Y = 9 else
"000000000000" when X = 252 AND Y = 9 else
"000000000000" when X = 253 AND Y = 9 else
"000000000000" when X = 254 AND Y = 9 else
"000000000000" when X = 255 AND Y = 9 else
"000000000000" when X = 256 AND Y = 9 else
"000000000000" when X = 257 AND Y = 9 else
"000000000000" when X = 258 AND Y = 9 else
"000000000000" when X = 259 AND Y = 9 else
"000000000000" when X = 260 AND Y = 9 else
"000000000000" when X = 261 AND Y = 9 else
"000000000000" when X = 262 AND Y = 9 else
"000000000000" when X = 263 AND Y = 9 else
"000000000000" when X = 264 AND Y = 9 else
"000000000000" when X = 265 AND Y = 9 else
"000000000000" when X = 266 AND Y = 9 else
"000000000000" when X = 267 AND Y = 9 else
"000000000000" when X = 268 AND Y = 9 else
"000000000000" when X = 269 AND Y = 9 else
"000000000000" when X = 270 AND Y = 9 else
"000000000000" when X = 271 AND Y = 9 else
"000000000000" when X = 272 AND Y = 9 else
"000000000000" when X = 273 AND Y = 9 else
"000000000000" when X = 274 AND Y = 9 else
"000000000000" when X = 275 AND Y = 9 else
"000000000000" when X = 276 AND Y = 9 else
"000000000000" when X = 277 AND Y = 9 else
"000000000000" when X = 278 AND Y = 9 else
"000000000000" when X = 279 AND Y = 9 else
"000000000000" when X = 280 AND Y = 9 else
"000000000000" when X = 281 AND Y = 9 else
"000000000000" when X = 282 AND Y = 9 else
"000000000000" when X = 283 AND Y = 9 else
"000000000000" when X = 284 AND Y = 9 else
"000000000000" when X = 285 AND Y = 9 else
"000000000000" when X = 286 AND Y = 9 else
"000000000000" when X = 287 AND Y = 9 else
"000000000000" when X = 288 AND Y = 9 else
"000000000000" when X = 289 AND Y = 9 else
"000000000000" when X = 290 AND Y = 9 else
"000000000000" when X = 291 AND Y = 9 else
"000000000000" when X = 292 AND Y = 9 else
"000000000000" when X = 293 AND Y = 9 else
"000000000000" when X = 294 AND Y = 9 else
"000000000000" when X = 295 AND Y = 9 else
"000000000000" when X = 296 AND Y = 9 else
"000000000000" when X = 297 AND Y = 9 else
"000000000000" when X = 298 AND Y = 9 else
"000000000000" when X = 299 AND Y = 9 else
"000000000000" when X = 300 AND Y = 9 else
"000000000000" when X = 301 AND Y = 9 else
"000000000000" when X = 302 AND Y = 9 else
"000000000000" when X = 303 AND Y = 9 else
"000000000000" when X = 304 AND Y = 9 else
"000000000000" when X = 305 AND Y = 9 else
"000000000000" when X = 306 AND Y = 9 else
"000000000000" when X = 307 AND Y = 9 else
"000000000000" when X = 308 AND Y = 9 else
"000000000000" when X = 309 AND Y = 9 else
"000000000000" when X = 310 AND Y = 9 else
"000000000000" when X = 311 AND Y = 9 else
"000000000000" when X = 312 AND Y = 9 else
"000000000000" when X = 313 AND Y = 9 else
"000000000000" when X = 314 AND Y = 9 else
"000000000000" when X = 315 AND Y = 9 else
"000000000000" when X = 316 AND Y = 9 else
"000000000000" when X = 317 AND Y = 9 else
"000000000000" when X = 318 AND Y = 9 else
"000000000000" when X = 319 AND Y = 9 else
"000000000000" when X = 320 AND Y = 9 else
"000000000000" when X = 321 AND Y = 9 else
"000000000000" when X = 322 AND Y = 9 else
"000000000000" when X = 323 AND Y = 9 else
"000000000000" when X = 324 AND Y = 9 else
"000000000000" when X = 0 AND Y = 10 else
"000000000000" when X = 1 AND Y = 10 else
"000000000000" when X = 2 AND Y = 10 else
"000000000000" when X = 3 AND Y = 10 else
"000000000000" when X = 4 AND Y = 10 else
"000000000000" when X = 5 AND Y = 10 else
"000000000000" when X = 6 AND Y = 10 else
"000000000000" when X = 7 AND Y = 10 else
"000000000000" when X = 8 AND Y = 10 else
"000000000000" when X = 9 AND Y = 10 else
"000000000000" when X = 10 AND Y = 10 else
"000000000000" when X = 11 AND Y = 10 else
"000000000000" when X = 12 AND Y = 10 else
"000000000000" when X = 13 AND Y = 10 else
"000000000000" when X = 14 AND Y = 10 else
"000000000000" when X = 15 AND Y = 10 else
"000000000000" when X = 16 AND Y = 10 else
"000000000000" when X = 17 AND Y = 10 else
"000000000000" when X = 18 AND Y = 10 else
"000000000000" when X = 19 AND Y = 10 else
"000000000000" when X = 20 AND Y = 10 else
"000000000000" when X = 21 AND Y = 10 else
"000000000000" when X = 22 AND Y = 10 else
"000000000000" when X = 23 AND Y = 10 else
"000000000000" when X = 24 AND Y = 10 else
"000000000000" when X = 25 AND Y = 10 else
"000000000000" when X = 26 AND Y = 10 else
"000000000000" when X = 27 AND Y = 10 else
"000000000000" when X = 28 AND Y = 10 else
"000000000000" when X = 29 AND Y = 10 else
"000000000000" when X = 30 AND Y = 10 else
"000000000000" when X = 31 AND Y = 10 else
"000000000000" when X = 32 AND Y = 10 else
"000000000000" when X = 33 AND Y = 10 else
"000000000000" when X = 34 AND Y = 10 else
"000000000000" when X = 35 AND Y = 10 else
"000000000000" when X = 36 AND Y = 10 else
"000000000000" when X = 37 AND Y = 10 else
"000000000000" when X = 38 AND Y = 10 else
"000000000000" when X = 39 AND Y = 10 else
"100010011101" when X = 40 AND Y = 10 else
"100010011101" when X = 41 AND Y = 10 else
"100010011101" when X = 42 AND Y = 10 else
"100010011101" when X = 43 AND Y = 10 else
"100010011101" when X = 44 AND Y = 10 else
"100010011101" when X = 45 AND Y = 10 else
"100010011101" when X = 46 AND Y = 10 else
"100010011101" when X = 47 AND Y = 10 else
"100010011101" when X = 48 AND Y = 10 else
"100010011101" when X = 49 AND Y = 10 else
"110111011111" when X = 50 AND Y = 10 else
"110111011111" when X = 51 AND Y = 10 else
"110111011111" when X = 52 AND Y = 10 else
"110111011111" when X = 53 AND Y = 10 else
"110111011111" when X = 54 AND Y = 10 else
"110111011111" when X = 55 AND Y = 10 else
"110111011111" when X = 56 AND Y = 10 else
"110111011111" when X = 57 AND Y = 10 else
"110111011111" when X = 58 AND Y = 10 else
"110111011111" when X = 59 AND Y = 10 else
"110111011111" when X = 60 AND Y = 10 else
"110111011111" when X = 61 AND Y = 10 else
"110111011111" when X = 62 AND Y = 10 else
"110111011111" when X = 63 AND Y = 10 else
"110111011111" when X = 64 AND Y = 10 else
"110111011111" when X = 65 AND Y = 10 else
"110111011111" when X = 66 AND Y = 10 else
"110111011111" when X = 67 AND Y = 10 else
"110111011111" when X = 68 AND Y = 10 else
"110111011111" when X = 69 AND Y = 10 else
"111111111111" when X = 70 AND Y = 10 else
"111111111111" when X = 71 AND Y = 10 else
"111111111111" when X = 72 AND Y = 10 else
"111111111111" when X = 73 AND Y = 10 else
"111111111111" when X = 74 AND Y = 10 else
"111111111111" when X = 75 AND Y = 10 else
"111111111111" when X = 76 AND Y = 10 else
"111111111111" when X = 77 AND Y = 10 else
"111111111111" when X = 78 AND Y = 10 else
"111111111111" when X = 79 AND Y = 10 else
"111111111111" when X = 80 AND Y = 10 else
"111111111111" when X = 81 AND Y = 10 else
"111111111111" when X = 82 AND Y = 10 else
"111111111111" when X = 83 AND Y = 10 else
"111111111111" when X = 84 AND Y = 10 else
"111111111111" when X = 85 AND Y = 10 else
"111111111111" when X = 86 AND Y = 10 else
"111111111111" when X = 87 AND Y = 10 else
"111111111111" when X = 88 AND Y = 10 else
"111111111111" when X = 89 AND Y = 10 else
"111111111111" when X = 90 AND Y = 10 else
"111111111111" when X = 91 AND Y = 10 else
"111111111111" when X = 92 AND Y = 10 else
"111111111111" when X = 93 AND Y = 10 else
"111111111111" when X = 94 AND Y = 10 else
"111111111111" when X = 95 AND Y = 10 else
"111111111111" when X = 96 AND Y = 10 else
"111111111111" when X = 97 AND Y = 10 else
"111111111111" when X = 98 AND Y = 10 else
"111111111111" when X = 99 AND Y = 10 else
"111111111111" when X = 100 AND Y = 10 else
"111111111111" when X = 101 AND Y = 10 else
"111111111111" when X = 102 AND Y = 10 else
"111111111111" when X = 103 AND Y = 10 else
"111111111111" when X = 104 AND Y = 10 else
"111111111111" when X = 105 AND Y = 10 else
"111111111111" when X = 106 AND Y = 10 else
"111111111111" when X = 107 AND Y = 10 else
"111111111111" when X = 108 AND Y = 10 else
"111111111111" when X = 109 AND Y = 10 else
"111111111111" when X = 110 AND Y = 10 else
"111111111111" when X = 111 AND Y = 10 else
"111111111111" when X = 112 AND Y = 10 else
"111111111111" when X = 113 AND Y = 10 else
"111111111111" when X = 114 AND Y = 10 else
"111111111111" when X = 115 AND Y = 10 else
"111111111111" when X = 116 AND Y = 10 else
"111111111111" when X = 117 AND Y = 10 else
"111111111111" when X = 118 AND Y = 10 else
"111111111111" when X = 119 AND Y = 10 else
"111111111111" when X = 120 AND Y = 10 else
"111111111111" when X = 121 AND Y = 10 else
"111111111111" when X = 122 AND Y = 10 else
"111111111111" when X = 123 AND Y = 10 else
"111111111111" when X = 124 AND Y = 10 else
"111111111111" when X = 125 AND Y = 10 else
"111111111111" when X = 126 AND Y = 10 else
"111111111111" when X = 127 AND Y = 10 else
"111111111111" when X = 128 AND Y = 10 else
"111111111111" when X = 129 AND Y = 10 else
"111111111111" when X = 130 AND Y = 10 else
"111111111111" when X = 131 AND Y = 10 else
"111111111111" when X = 132 AND Y = 10 else
"111111111111" when X = 133 AND Y = 10 else
"111111111111" when X = 134 AND Y = 10 else
"111111111111" when X = 135 AND Y = 10 else
"111111111111" when X = 136 AND Y = 10 else
"111111111111" when X = 137 AND Y = 10 else
"111111111111" when X = 138 AND Y = 10 else
"111111111111" when X = 139 AND Y = 10 else
"111111111111" when X = 140 AND Y = 10 else
"111111111111" when X = 141 AND Y = 10 else
"111111111111" when X = 142 AND Y = 10 else
"111111111111" when X = 143 AND Y = 10 else
"111111111111" when X = 144 AND Y = 10 else
"111111111111" when X = 145 AND Y = 10 else
"111111111111" when X = 146 AND Y = 10 else
"111111111111" when X = 147 AND Y = 10 else
"111111111111" when X = 148 AND Y = 10 else
"111111111111" when X = 149 AND Y = 10 else
"000000000000" when X = 150 AND Y = 10 else
"000000000000" when X = 151 AND Y = 10 else
"000000000000" when X = 152 AND Y = 10 else
"000000000000" when X = 153 AND Y = 10 else
"000000000000" when X = 154 AND Y = 10 else
"000000000000" when X = 155 AND Y = 10 else
"000000000000" when X = 156 AND Y = 10 else
"000000000000" when X = 157 AND Y = 10 else
"000000000000" when X = 158 AND Y = 10 else
"000000000000" when X = 159 AND Y = 10 else
"000000000000" when X = 160 AND Y = 10 else
"000000000000" when X = 161 AND Y = 10 else
"000000000000" when X = 162 AND Y = 10 else
"000000000000" when X = 163 AND Y = 10 else
"000000000000" when X = 164 AND Y = 10 else
"000000000000" when X = 165 AND Y = 10 else
"000000000000" when X = 166 AND Y = 10 else
"000000000000" when X = 167 AND Y = 10 else
"000000000000" when X = 168 AND Y = 10 else
"000000000000" when X = 169 AND Y = 10 else
"000000000000" when X = 170 AND Y = 10 else
"000000000000" when X = 171 AND Y = 10 else
"000000000000" when X = 172 AND Y = 10 else
"000000000000" when X = 173 AND Y = 10 else
"000000000000" when X = 174 AND Y = 10 else
"000000000000" when X = 175 AND Y = 10 else
"000000000000" when X = 176 AND Y = 10 else
"000000000000" when X = 177 AND Y = 10 else
"000000000000" when X = 178 AND Y = 10 else
"000000000000" when X = 179 AND Y = 10 else
"000000000000" when X = 180 AND Y = 10 else
"000000000000" when X = 181 AND Y = 10 else
"000000000000" when X = 182 AND Y = 10 else
"000000000000" when X = 183 AND Y = 10 else
"000000000000" when X = 184 AND Y = 10 else
"000000000000" when X = 185 AND Y = 10 else
"000000000000" when X = 186 AND Y = 10 else
"000000000000" when X = 187 AND Y = 10 else
"000000000000" when X = 188 AND Y = 10 else
"000000000000" when X = 189 AND Y = 10 else
"000000000000" when X = 190 AND Y = 10 else
"000000000000" when X = 191 AND Y = 10 else
"000000000000" when X = 192 AND Y = 10 else
"000000000000" when X = 193 AND Y = 10 else
"000000000000" when X = 194 AND Y = 10 else
"000000000000" when X = 195 AND Y = 10 else
"000000000000" when X = 196 AND Y = 10 else
"000000000000" when X = 197 AND Y = 10 else
"000000000000" when X = 198 AND Y = 10 else
"000000000000" when X = 199 AND Y = 10 else
"000000000000" when X = 200 AND Y = 10 else
"000000000000" when X = 201 AND Y = 10 else
"000000000000" when X = 202 AND Y = 10 else
"000000000000" when X = 203 AND Y = 10 else
"000000000000" when X = 204 AND Y = 10 else
"000000000000" when X = 205 AND Y = 10 else
"000000000000" when X = 206 AND Y = 10 else
"000000000000" when X = 207 AND Y = 10 else
"000000000000" when X = 208 AND Y = 10 else
"000000000000" when X = 209 AND Y = 10 else
"000000000000" when X = 210 AND Y = 10 else
"000000000000" when X = 211 AND Y = 10 else
"000000000000" when X = 212 AND Y = 10 else
"000000000000" when X = 213 AND Y = 10 else
"000000000000" when X = 214 AND Y = 10 else
"000000000000" when X = 215 AND Y = 10 else
"000000000000" when X = 216 AND Y = 10 else
"000000000000" when X = 217 AND Y = 10 else
"000000000000" when X = 218 AND Y = 10 else
"000000000000" when X = 219 AND Y = 10 else
"000000000000" when X = 220 AND Y = 10 else
"000000000000" when X = 221 AND Y = 10 else
"000000000000" when X = 222 AND Y = 10 else
"000000000000" when X = 223 AND Y = 10 else
"000000000000" when X = 224 AND Y = 10 else
"000000000000" when X = 225 AND Y = 10 else
"000000000000" when X = 226 AND Y = 10 else
"000000000000" when X = 227 AND Y = 10 else
"000000000000" when X = 228 AND Y = 10 else
"000000000000" when X = 229 AND Y = 10 else
"000000000000" when X = 230 AND Y = 10 else
"000000000000" when X = 231 AND Y = 10 else
"000000000000" when X = 232 AND Y = 10 else
"000000000000" when X = 233 AND Y = 10 else
"000000000000" when X = 234 AND Y = 10 else
"000000000000" when X = 235 AND Y = 10 else
"000000000000" when X = 236 AND Y = 10 else
"000000000000" when X = 237 AND Y = 10 else
"000000000000" when X = 238 AND Y = 10 else
"000000000000" when X = 239 AND Y = 10 else
"000000000000" when X = 240 AND Y = 10 else
"000000000000" when X = 241 AND Y = 10 else
"000000000000" when X = 242 AND Y = 10 else
"000000000000" when X = 243 AND Y = 10 else
"000000000000" when X = 244 AND Y = 10 else
"000000000000" when X = 245 AND Y = 10 else
"000000000000" when X = 246 AND Y = 10 else
"000000000000" when X = 247 AND Y = 10 else
"000000000000" when X = 248 AND Y = 10 else
"000000000000" when X = 249 AND Y = 10 else
"000000000000" when X = 250 AND Y = 10 else
"000000000000" when X = 251 AND Y = 10 else
"000000000000" when X = 252 AND Y = 10 else
"000000000000" when X = 253 AND Y = 10 else
"000000000000" when X = 254 AND Y = 10 else
"000000000000" when X = 255 AND Y = 10 else
"000000000000" when X = 256 AND Y = 10 else
"000000000000" when X = 257 AND Y = 10 else
"000000000000" when X = 258 AND Y = 10 else
"000000000000" when X = 259 AND Y = 10 else
"000000000000" when X = 260 AND Y = 10 else
"000000000000" when X = 261 AND Y = 10 else
"000000000000" when X = 262 AND Y = 10 else
"000000000000" when X = 263 AND Y = 10 else
"000000000000" when X = 264 AND Y = 10 else
"000000000000" when X = 265 AND Y = 10 else
"000000000000" when X = 266 AND Y = 10 else
"000000000000" when X = 267 AND Y = 10 else
"000000000000" when X = 268 AND Y = 10 else
"000000000000" when X = 269 AND Y = 10 else
"000000000000" when X = 270 AND Y = 10 else
"000000000000" when X = 271 AND Y = 10 else
"000000000000" when X = 272 AND Y = 10 else
"000000000000" when X = 273 AND Y = 10 else
"000000000000" when X = 274 AND Y = 10 else
"000000000000" when X = 275 AND Y = 10 else
"000000000000" when X = 276 AND Y = 10 else
"000000000000" when X = 277 AND Y = 10 else
"000000000000" when X = 278 AND Y = 10 else
"000000000000" when X = 279 AND Y = 10 else
"000000000000" when X = 280 AND Y = 10 else
"000000000000" when X = 281 AND Y = 10 else
"000000000000" when X = 282 AND Y = 10 else
"000000000000" when X = 283 AND Y = 10 else
"000000000000" when X = 284 AND Y = 10 else
"000000000000" when X = 285 AND Y = 10 else
"000000000000" when X = 286 AND Y = 10 else
"000000000000" when X = 287 AND Y = 10 else
"000000000000" when X = 288 AND Y = 10 else
"000000000000" when X = 289 AND Y = 10 else
"000000000000" when X = 290 AND Y = 10 else
"000000000000" when X = 291 AND Y = 10 else
"000000000000" when X = 292 AND Y = 10 else
"000000000000" when X = 293 AND Y = 10 else
"000000000000" when X = 294 AND Y = 10 else
"000000000000" when X = 295 AND Y = 10 else
"000000000000" when X = 296 AND Y = 10 else
"000000000000" when X = 297 AND Y = 10 else
"000000000000" when X = 298 AND Y = 10 else
"000000000000" when X = 299 AND Y = 10 else
"000000000000" when X = 300 AND Y = 10 else
"000000000000" when X = 301 AND Y = 10 else
"000000000000" when X = 302 AND Y = 10 else
"000000000000" when X = 303 AND Y = 10 else
"000000000000" when X = 304 AND Y = 10 else
"000000000000" when X = 305 AND Y = 10 else
"000000000000" when X = 306 AND Y = 10 else
"000000000000" when X = 307 AND Y = 10 else
"000000000000" when X = 308 AND Y = 10 else
"000000000000" when X = 309 AND Y = 10 else
"000000000000" when X = 310 AND Y = 10 else
"000000000000" when X = 311 AND Y = 10 else
"000000000000" when X = 312 AND Y = 10 else
"000000000000" when X = 313 AND Y = 10 else
"000000000000" when X = 314 AND Y = 10 else
"000000000000" when X = 315 AND Y = 10 else
"000000000000" when X = 316 AND Y = 10 else
"000000000000" when X = 317 AND Y = 10 else
"000000000000" when X = 318 AND Y = 10 else
"000000000000" when X = 319 AND Y = 10 else
"000000000000" when X = 320 AND Y = 10 else
"000000000000" when X = 321 AND Y = 10 else
"000000000000" when X = 322 AND Y = 10 else
"000000000000" when X = 323 AND Y = 10 else
"000000000000" when X = 324 AND Y = 10 else
"000000000000" when X = 0 AND Y = 11 else
"000000000000" when X = 1 AND Y = 11 else
"000000000000" when X = 2 AND Y = 11 else
"000000000000" when X = 3 AND Y = 11 else
"000000000000" when X = 4 AND Y = 11 else
"000000000000" when X = 5 AND Y = 11 else
"000000000000" when X = 6 AND Y = 11 else
"000000000000" when X = 7 AND Y = 11 else
"000000000000" when X = 8 AND Y = 11 else
"000000000000" when X = 9 AND Y = 11 else
"000000000000" when X = 10 AND Y = 11 else
"000000000000" when X = 11 AND Y = 11 else
"000000000000" when X = 12 AND Y = 11 else
"000000000000" when X = 13 AND Y = 11 else
"000000000000" when X = 14 AND Y = 11 else
"000000000000" when X = 15 AND Y = 11 else
"000000000000" when X = 16 AND Y = 11 else
"000000000000" when X = 17 AND Y = 11 else
"000000000000" when X = 18 AND Y = 11 else
"000000000000" when X = 19 AND Y = 11 else
"000000000000" when X = 20 AND Y = 11 else
"000000000000" when X = 21 AND Y = 11 else
"000000000000" when X = 22 AND Y = 11 else
"000000000000" when X = 23 AND Y = 11 else
"000000000000" when X = 24 AND Y = 11 else
"000000000000" when X = 25 AND Y = 11 else
"000000000000" when X = 26 AND Y = 11 else
"000000000000" when X = 27 AND Y = 11 else
"000000000000" when X = 28 AND Y = 11 else
"000000000000" when X = 29 AND Y = 11 else
"000000000000" when X = 30 AND Y = 11 else
"000000000000" when X = 31 AND Y = 11 else
"000000000000" when X = 32 AND Y = 11 else
"000000000000" when X = 33 AND Y = 11 else
"000000000000" when X = 34 AND Y = 11 else
"000000000000" when X = 35 AND Y = 11 else
"000000000000" when X = 36 AND Y = 11 else
"000000000000" when X = 37 AND Y = 11 else
"000000000000" when X = 38 AND Y = 11 else
"000000000000" when X = 39 AND Y = 11 else
"100010011101" when X = 40 AND Y = 11 else
"100010011101" when X = 41 AND Y = 11 else
"100010011101" when X = 42 AND Y = 11 else
"100010011101" when X = 43 AND Y = 11 else
"100010011101" when X = 44 AND Y = 11 else
"100010011101" when X = 45 AND Y = 11 else
"100010011101" when X = 46 AND Y = 11 else
"100010011101" when X = 47 AND Y = 11 else
"100010011101" when X = 48 AND Y = 11 else
"100010011101" when X = 49 AND Y = 11 else
"110111011111" when X = 50 AND Y = 11 else
"110111011111" when X = 51 AND Y = 11 else
"110111011111" when X = 52 AND Y = 11 else
"110111011111" when X = 53 AND Y = 11 else
"110111011111" when X = 54 AND Y = 11 else
"110111011111" when X = 55 AND Y = 11 else
"110111011111" when X = 56 AND Y = 11 else
"110111011111" when X = 57 AND Y = 11 else
"110111011111" when X = 58 AND Y = 11 else
"110111011111" when X = 59 AND Y = 11 else
"110111011111" when X = 60 AND Y = 11 else
"110111011111" when X = 61 AND Y = 11 else
"110111011111" when X = 62 AND Y = 11 else
"110111011111" when X = 63 AND Y = 11 else
"110111011111" when X = 64 AND Y = 11 else
"110111011111" when X = 65 AND Y = 11 else
"110111011111" when X = 66 AND Y = 11 else
"110111011111" when X = 67 AND Y = 11 else
"110111011111" when X = 68 AND Y = 11 else
"110111011111" when X = 69 AND Y = 11 else
"111111111111" when X = 70 AND Y = 11 else
"111111111111" when X = 71 AND Y = 11 else
"111111111111" when X = 72 AND Y = 11 else
"111111111111" when X = 73 AND Y = 11 else
"111111111111" when X = 74 AND Y = 11 else
"111111111111" when X = 75 AND Y = 11 else
"111111111111" when X = 76 AND Y = 11 else
"111111111111" when X = 77 AND Y = 11 else
"111111111111" when X = 78 AND Y = 11 else
"111111111111" when X = 79 AND Y = 11 else
"111111111111" when X = 80 AND Y = 11 else
"111111111111" when X = 81 AND Y = 11 else
"111111111111" when X = 82 AND Y = 11 else
"111111111111" when X = 83 AND Y = 11 else
"111111111111" when X = 84 AND Y = 11 else
"111111111111" when X = 85 AND Y = 11 else
"111111111111" when X = 86 AND Y = 11 else
"111111111111" when X = 87 AND Y = 11 else
"111111111111" when X = 88 AND Y = 11 else
"111111111111" when X = 89 AND Y = 11 else
"111111111111" when X = 90 AND Y = 11 else
"111111111111" when X = 91 AND Y = 11 else
"111111111111" when X = 92 AND Y = 11 else
"111111111111" when X = 93 AND Y = 11 else
"111111111111" when X = 94 AND Y = 11 else
"111111111111" when X = 95 AND Y = 11 else
"111111111111" when X = 96 AND Y = 11 else
"111111111111" when X = 97 AND Y = 11 else
"111111111111" when X = 98 AND Y = 11 else
"111111111111" when X = 99 AND Y = 11 else
"111111111111" when X = 100 AND Y = 11 else
"111111111111" when X = 101 AND Y = 11 else
"111111111111" when X = 102 AND Y = 11 else
"111111111111" when X = 103 AND Y = 11 else
"111111111111" when X = 104 AND Y = 11 else
"111111111111" when X = 105 AND Y = 11 else
"111111111111" when X = 106 AND Y = 11 else
"111111111111" when X = 107 AND Y = 11 else
"111111111111" when X = 108 AND Y = 11 else
"111111111111" when X = 109 AND Y = 11 else
"111111111111" when X = 110 AND Y = 11 else
"111111111111" when X = 111 AND Y = 11 else
"111111111111" when X = 112 AND Y = 11 else
"111111111111" when X = 113 AND Y = 11 else
"111111111111" when X = 114 AND Y = 11 else
"111111111111" when X = 115 AND Y = 11 else
"111111111111" when X = 116 AND Y = 11 else
"111111111111" when X = 117 AND Y = 11 else
"111111111111" when X = 118 AND Y = 11 else
"111111111111" when X = 119 AND Y = 11 else
"111111111111" when X = 120 AND Y = 11 else
"111111111111" when X = 121 AND Y = 11 else
"111111111111" when X = 122 AND Y = 11 else
"111111111111" when X = 123 AND Y = 11 else
"111111111111" when X = 124 AND Y = 11 else
"111111111111" when X = 125 AND Y = 11 else
"111111111111" when X = 126 AND Y = 11 else
"111111111111" when X = 127 AND Y = 11 else
"111111111111" when X = 128 AND Y = 11 else
"111111111111" when X = 129 AND Y = 11 else
"111111111111" when X = 130 AND Y = 11 else
"111111111111" when X = 131 AND Y = 11 else
"111111111111" when X = 132 AND Y = 11 else
"111111111111" when X = 133 AND Y = 11 else
"111111111111" when X = 134 AND Y = 11 else
"111111111111" when X = 135 AND Y = 11 else
"111111111111" when X = 136 AND Y = 11 else
"111111111111" when X = 137 AND Y = 11 else
"111111111111" when X = 138 AND Y = 11 else
"111111111111" when X = 139 AND Y = 11 else
"111111111111" when X = 140 AND Y = 11 else
"111111111111" when X = 141 AND Y = 11 else
"111111111111" when X = 142 AND Y = 11 else
"111111111111" when X = 143 AND Y = 11 else
"111111111111" when X = 144 AND Y = 11 else
"111111111111" when X = 145 AND Y = 11 else
"111111111111" when X = 146 AND Y = 11 else
"111111111111" when X = 147 AND Y = 11 else
"111111111111" when X = 148 AND Y = 11 else
"111111111111" when X = 149 AND Y = 11 else
"000000000000" when X = 150 AND Y = 11 else
"000000000000" when X = 151 AND Y = 11 else
"000000000000" when X = 152 AND Y = 11 else
"000000000000" when X = 153 AND Y = 11 else
"000000000000" when X = 154 AND Y = 11 else
"000000000000" when X = 155 AND Y = 11 else
"000000000000" when X = 156 AND Y = 11 else
"000000000000" when X = 157 AND Y = 11 else
"000000000000" when X = 158 AND Y = 11 else
"000000000000" when X = 159 AND Y = 11 else
"000000000000" when X = 160 AND Y = 11 else
"000000000000" when X = 161 AND Y = 11 else
"000000000000" when X = 162 AND Y = 11 else
"000000000000" when X = 163 AND Y = 11 else
"000000000000" when X = 164 AND Y = 11 else
"000000000000" when X = 165 AND Y = 11 else
"000000000000" when X = 166 AND Y = 11 else
"000000000000" when X = 167 AND Y = 11 else
"000000000000" when X = 168 AND Y = 11 else
"000000000000" when X = 169 AND Y = 11 else
"000000000000" when X = 170 AND Y = 11 else
"000000000000" when X = 171 AND Y = 11 else
"000000000000" when X = 172 AND Y = 11 else
"000000000000" when X = 173 AND Y = 11 else
"000000000000" when X = 174 AND Y = 11 else
"000000000000" when X = 175 AND Y = 11 else
"000000000000" when X = 176 AND Y = 11 else
"000000000000" when X = 177 AND Y = 11 else
"000000000000" when X = 178 AND Y = 11 else
"000000000000" when X = 179 AND Y = 11 else
"000000000000" when X = 180 AND Y = 11 else
"000000000000" when X = 181 AND Y = 11 else
"000000000000" when X = 182 AND Y = 11 else
"000000000000" when X = 183 AND Y = 11 else
"000000000000" when X = 184 AND Y = 11 else
"000000000000" when X = 185 AND Y = 11 else
"000000000000" when X = 186 AND Y = 11 else
"000000000000" when X = 187 AND Y = 11 else
"000000000000" when X = 188 AND Y = 11 else
"000000000000" when X = 189 AND Y = 11 else
"000000000000" when X = 190 AND Y = 11 else
"000000000000" when X = 191 AND Y = 11 else
"000000000000" when X = 192 AND Y = 11 else
"000000000000" when X = 193 AND Y = 11 else
"000000000000" when X = 194 AND Y = 11 else
"000000000000" when X = 195 AND Y = 11 else
"000000000000" when X = 196 AND Y = 11 else
"000000000000" when X = 197 AND Y = 11 else
"000000000000" when X = 198 AND Y = 11 else
"000000000000" when X = 199 AND Y = 11 else
"000000000000" when X = 200 AND Y = 11 else
"000000000000" when X = 201 AND Y = 11 else
"000000000000" when X = 202 AND Y = 11 else
"000000000000" when X = 203 AND Y = 11 else
"000000000000" when X = 204 AND Y = 11 else
"000000000000" when X = 205 AND Y = 11 else
"000000000000" when X = 206 AND Y = 11 else
"000000000000" when X = 207 AND Y = 11 else
"000000000000" when X = 208 AND Y = 11 else
"000000000000" when X = 209 AND Y = 11 else
"000000000000" when X = 210 AND Y = 11 else
"000000000000" when X = 211 AND Y = 11 else
"000000000000" when X = 212 AND Y = 11 else
"000000000000" when X = 213 AND Y = 11 else
"000000000000" when X = 214 AND Y = 11 else
"000000000000" when X = 215 AND Y = 11 else
"000000000000" when X = 216 AND Y = 11 else
"000000000000" when X = 217 AND Y = 11 else
"000000000000" when X = 218 AND Y = 11 else
"000000000000" when X = 219 AND Y = 11 else
"000000000000" when X = 220 AND Y = 11 else
"000000000000" when X = 221 AND Y = 11 else
"000000000000" when X = 222 AND Y = 11 else
"000000000000" when X = 223 AND Y = 11 else
"000000000000" when X = 224 AND Y = 11 else
"000000000000" when X = 225 AND Y = 11 else
"000000000000" when X = 226 AND Y = 11 else
"000000000000" when X = 227 AND Y = 11 else
"000000000000" when X = 228 AND Y = 11 else
"000000000000" when X = 229 AND Y = 11 else
"000000000000" when X = 230 AND Y = 11 else
"000000000000" when X = 231 AND Y = 11 else
"000000000000" when X = 232 AND Y = 11 else
"000000000000" when X = 233 AND Y = 11 else
"000000000000" when X = 234 AND Y = 11 else
"000000000000" when X = 235 AND Y = 11 else
"000000000000" when X = 236 AND Y = 11 else
"000000000000" when X = 237 AND Y = 11 else
"000000000000" when X = 238 AND Y = 11 else
"000000000000" when X = 239 AND Y = 11 else
"000000000000" when X = 240 AND Y = 11 else
"000000000000" when X = 241 AND Y = 11 else
"000000000000" when X = 242 AND Y = 11 else
"000000000000" when X = 243 AND Y = 11 else
"000000000000" when X = 244 AND Y = 11 else
"000000000000" when X = 245 AND Y = 11 else
"000000000000" when X = 246 AND Y = 11 else
"000000000000" when X = 247 AND Y = 11 else
"000000000000" when X = 248 AND Y = 11 else
"000000000000" when X = 249 AND Y = 11 else
"000000000000" when X = 250 AND Y = 11 else
"000000000000" when X = 251 AND Y = 11 else
"000000000000" when X = 252 AND Y = 11 else
"000000000000" when X = 253 AND Y = 11 else
"000000000000" when X = 254 AND Y = 11 else
"000000000000" when X = 255 AND Y = 11 else
"000000000000" when X = 256 AND Y = 11 else
"000000000000" when X = 257 AND Y = 11 else
"000000000000" when X = 258 AND Y = 11 else
"000000000000" when X = 259 AND Y = 11 else
"000000000000" when X = 260 AND Y = 11 else
"000000000000" when X = 261 AND Y = 11 else
"000000000000" when X = 262 AND Y = 11 else
"000000000000" when X = 263 AND Y = 11 else
"000000000000" when X = 264 AND Y = 11 else
"000000000000" when X = 265 AND Y = 11 else
"000000000000" when X = 266 AND Y = 11 else
"000000000000" when X = 267 AND Y = 11 else
"000000000000" when X = 268 AND Y = 11 else
"000000000000" when X = 269 AND Y = 11 else
"000000000000" when X = 270 AND Y = 11 else
"000000000000" when X = 271 AND Y = 11 else
"000000000000" when X = 272 AND Y = 11 else
"000000000000" when X = 273 AND Y = 11 else
"000000000000" when X = 274 AND Y = 11 else
"000000000000" when X = 275 AND Y = 11 else
"000000000000" when X = 276 AND Y = 11 else
"000000000000" when X = 277 AND Y = 11 else
"000000000000" when X = 278 AND Y = 11 else
"000000000000" when X = 279 AND Y = 11 else
"000000000000" when X = 280 AND Y = 11 else
"000000000000" when X = 281 AND Y = 11 else
"000000000000" when X = 282 AND Y = 11 else
"000000000000" when X = 283 AND Y = 11 else
"000000000000" when X = 284 AND Y = 11 else
"000000000000" when X = 285 AND Y = 11 else
"000000000000" when X = 286 AND Y = 11 else
"000000000000" when X = 287 AND Y = 11 else
"000000000000" when X = 288 AND Y = 11 else
"000000000000" when X = 289 AND Y = 11 else
"000000000000" when X = 290 AND Y = 11 else
"000000000000" when X = 291 AND Y = 11 else
"000000000000" when X = 292 AND Y = 11 else
"000000000000" when X = 293 AND Y = 11 else
"000000000000" when X = 294 AND Y = 11 else
"000000000000" when X = 295 AND Y = 11 else
"000000000000" when X = 296 AND Y = 11 else
"000000000000" when X = 297 AND Y = 11 else
"000000000000" when X = 298 AND Y = 11 else
"000000000000" when X = 299 AND Y = 11 else
"000000000000" when X = 300 AND Y = 11 else
"000000000000" when X = 301 AND Y = 11 else
"000000000000" when X = 302 AND Y = 11 else
"000000000000" when X = 303 AND Y = 11 else
"000000000000" when X = 304 AND Y = 11 else
"000000000000" when X = 305 AND Y = 11 else
"000000000000" when X = 306 AND Y = 11 else
"000000000000" when X = 307 AND Y = 11 else
"000000000000" when X = 308 AND Y = 11 else
"000000000000" when X = 309 AND Y = 11 else
"000000000000" when X = 310 AND Y = 11 else
"000000000000" when X = 311 AND Y = 11 else
"000000000000" when X = 312 AND Y = 11 else
"000000000000" when X = 313 AND Y = 11 else
"000000000000" when X = 314 AND Y = 11 else
"000000000000" when X = 315 AND Y = 11 else
"000000000000" when X = 316 AND Y = 11 else
"000000000000" when X = 317 AND Y = 11 else
"000000000000" when X = 318 AND Y = 11 else
"000000000000" when X = 319 AND Y = 11 else
"000000000000" when X = 320 AND Y = 11 else
"000000000000" when X = 321 AND Y = 11 else
"000000000000" when X = 322 AND Y = 11 else
"000000000000" when X = 323 AND Y = 11 else
"000000000000" when X = 324 AND Y = 11 else
"000000000000" when X = 0 AND Y = 12 else
"000000000000" when X = 1 AND Y = 12 else
"000000000000" when X = 2 AND Y = 12 else
"000000000000" when X = 3 AND Y = 12 else
"000000000000" when X = 4 AND Y = 12 else
"000000000000" when X = 5 AND Y = 12 else
"000000000000" when X = 6 AND Y = 12 else
"000000000000" when X = 7 AND Y = 12 else
"000000000000" when X = 8 AND Y = 12 else
"000000000000" when X = 9 AND Y = 12 else
"000000000000" when X = 10 AND Y = 12 else
"000000000000" when X = 11 AND Y = 12 else
"000000000000" when X = 12 AND Y = 12 else
"000000000000" when X = 13 AND Y = 12 else
"000000000000" when X = 14 AND Y = 12 else
"000000000000" when X = 15 AND Y = 12 else
"000000000000" when X = 16 AND Y = 12 else
"000000000000" when X = 17 AND Y = 12 else
"000000000000" when X = 18 AND Y = 12 else
"000000000000" when X = 19 AND Y = 12 else
"000000000000" when X = 20 AND Y = 12 else
"000000000000" when X = 21 AND Y = 12 else
"000000000000" when X = 22 AND Y = 12 else
"000000000000" when X = 23 AND Y = 12 else
"000000000000" when X = 24 AND Y = 12 else
"000000000000" when X = 25 AND Y = 12 else
"000000000000" when X = 26 AND Y = 12 else
"000000000000" when X = 27 AND Y = 12 else
"000000000000" when X = 28 AND Y = 12 else
"000000000000" when X = 29 AND Y = 12 else
"000000000000" when X = 30 AND Y = 12 else
"000000000000" when X = 31 AND Y = 12 else
"000000000000" when X = 32 AND Y = 12 else
"000000000000" when X = 33 AND Y = 12 else
"000000000000" when X = 34 AND Y = 12 else
"000000000000" when X = 35 AND Y = 12 else
"000000000000" when X = 36 AND Y = 12 else
"000000000000" when X = 37 AND Y = 12 else
"000000000000" when X = 38 AND Y = 12 else
"000000000000" when X = 39 AND Y = 12 else
"100010011101" when X = 40 AND Y = 12 else
"100010011101" when X = 41 AND Y = 12 else
"100010011101" when X = 42 AND Y = 12 else
"100010011101" when X = 43 AND Y = 12 else
"100010011101" when X = 44 AND Y = 12 else
"100010011101" when X = 45 AND Y = 12 else
"100010011101" when X = 46 AND Y = 12 else
"100010011101" when X = 47 AND Y = 12 else
"100010011101" when X = 48 AND Y = 12 else
"100010011101" when X = 49 AND Y = 12 else
"110111011111" when X = 50 AND Y = 12 else
"110111011111" when X = 51 AND Y = 12 else
"110111011111" when X = 52 AND Y = 12 else
"110111011111" when X = 53 AND Y = 12 else
"110111011111" when X = 54 AND Y = 12 else
"110111011111" when X = 55 AND Y = 12 else
"110111011111" when X = 56 AND Y = 12 else
"110111011111" when X = 57 AND Y = 12 else
"110111011111" when X = 58 AND Y = 12 else
"110111011111" when X = 59 AND Y = 12 else
"110111011111" when X = 60 AND Y = 12 else
"110111011111" when X = 61 AND Y = 12 else
"110111011111" when X = 62 AND Y = 12 else
"110111011111" when X = 63 AND Y = 12 else
"110111011111" when X = 64 AND Y = 12 else
"110111011111" when X = 65 AND Y = 12 else
"110111011111" when X = 66 AND Y = 12 else
"110111011111" when X = 67 AND Y = 12 else
"110111011111" when X = 68 AND Y = 12 else
"110111011111" when X = 69 AND Y = 12 else
"111111111111" when X = 70 AND Y = 12 else
"111111111111" when X = 71 AND Y = 12 else
"111111111111" when X = 72 AND Y = 12 else
"111111111111" when X = 73 AND Y = 12 else
"111111111111" when X = 74 AND Y = 12 else
"111111111111" when X = 75 AND Y = 12 else
"111111111111" when X = 76 AND Y = 12 else
"111111111111" when X = 77 AND Y = 12 else
"111111111111" when X = 78 AND Y = 12 else
"111111111111" when X = 79 AND Y = 12 else
"111111111111" when X = 80 AND Y = 12 else
"111111111111" when X = 81 AND Y = 12 else
"111111111111" when X = 82 AND Y = 12 else
"111111111111" when X = 83 AND Y = 12 else
"111111111111" when X = 84 AND Y = 12 else
"111111111111" when X = 85 AND Y = 12 else
"111111111111" when X = 86 AND Y = 12 else
"111111111111" when X = 87 AND Y = 12 else
"111111111111" when X = 88 AND Y = 12 else
"111111111111" when X = 89 AND Y = 12 else
"111111111111" when X = 90 AND Y = 12 else
"111111111111" when X = 91 AND Y = 12 else
"111111111111" when X = 92 AND Y = 12 else
"111111111111" when X = 93 AND Y = 12 else
"111111111111" when X = 94 AND Y = 12 else
"111111111111" when X = 95 AND Y = 12 else
"111111111111" when X = 96 AND Y = 12 else
"111111111111" when X = 97 AND Y = 12 else
"111111111111" when X = 98 AND Y = 12 else
"111111111111" when X = 99 AND Y = 12 else
"111111111111" when X = 100 AND Y = 12 else
"111111111111" when X = 101 AND Y = 12 else
"111111111111" when X = 102 AND Y = 12 else
"111111111111" when X = 103 AND Y = 12 else
"111111111111" when X = 104 AND Y = 12 else
"111111111111" when X = 105 AND Y = 12 else
"111111111111" when X = 106 AND Y = 12 else
"111111111111" when X = 107 AND Y = 12 else
"111111111111" when X = 108 AND Y = 12 else
"111111111111" when X = 109 AND Y = 12 else
"111111111111" when X = 110 AND Y = 12 else
"111111111111" when X = 111 AND Y = 12 else
"111111111111" when X = 112 AND Y = 12 else
"111111111111" when X = 113 AND Y = 12 else
"111111111111" when X = 114 AND Y = 12 else
"111111111111" when X = 115 AND Y = 12 else
"111111111111" when X = 116 AND Y = 12 else
"111111111111" when X = 117 AND Y = 12 else
"111111111111" when X = 118 AND Y = 12 else
"111111111111" when X = 119 AND Y = 12 else
"111111111111" when X = 120 AND Y = 12 else
"111111111111" when X = 121 AND Y = 12 else
"111111111111" when X = 122 AND Y = 12 else
"111111111111" when X = 123 AND Y = 12 else
"111111111111" when X = 124 AND Y = 12 else
"111111111111" when X = 125 AND Y = 12 else
"111111111111" when X = 126 AND Y = 12 else
"111111111111" when X = 127 AND Y = 12 else
"111111111111" when X = 128 AND Y = 12 else
"111111111111" when X = 129 AND Y = 12 else
"111111111111" when X = 130 AND Y = 12 else
"111111111111" when X = 131 AND Y = 12 else
"111111111111" when X = 132 AND Y = 12 else
"111111111111" when X = 133 AND Y = 12 else
"111111111111" when X = 134 AND Y = 12 else
"111111111111" when X = 135 AND Y = 12 else
"111111111111" when X = 136 AND Y = 12 else
"111111111111" when X = 137 AND Y = 12 else
"111111111111" when X = 138 AND Y = 12 else
"111111111111" when X = 139 AND Y = 12 else
"111111111111" when X = 140 AND Y = 12 else
"111111111111" when X = 141 AND Y = 12 else
"111111111111" when X = 142 AND Y = 12 else
"111111111111" when X = 143 AND Y = 12 else
"111111111111" when X = 144 AND Y = 12 else
"111111111111" when X = 145 AND Y = 12 else
"111111111111" when X = 146 AND Y = 12 else
"111111111111" when X = 147 AND Y = 12 else
"111111111111" when X = 148 AND Y = 12 else
"111111111111" when X = 149 AND Y = 12 else
"000000000000" when X = 150 AND Y = 12 else
"000000000000" when X = 151 AND Y = 12 else
"000000000000" when X = 152 AND Y = 12 else
"000000000000" when X = 153 AND Y = 12 else
"000000000000" when X = 154 AND Y = 12 else
"000000000000" when X = 155 AND Y = 12 else
"000000000000" when X = 156 AND Y = 12 else
"000000000000" when X = 157 AND Y = 12 else
"000000000000" when X = 158 AND Y = 12 else
"000000000000" when X = 159 AND Y = 12 else
"000000000000" when X = 160 AND Y = 12 else
"000000000000" when X = 161 AND Y = 12 else
"000000000000" when X = 162 AND Y = 12 else
"000000000000" when X = 163 AND Y = 12 else
"000000000000" when X = 164 AND Y = 12 else
"000000000000" when X = 165 AND Y = 12 else
"000000000000" when X = 166 AND Y = 12 else
"000000000000" when X = 167 AND Y = 12 else
"000000000000" when X = 168 AND Y = 12 else
"000000000000" when X = 169 AND Y = 12 else
"000000000000" when X = 170 AND Y = 12 else
"000000000000" when X = 171 AND Y = 12 else
"000000000000" when X = 172 AND Y = 12 else
"000000000000" when X = 173 AND Y = 12 else
"000000000000" when X = 174 AND Y = 12 else
"000000000000" when X = 175 AND Y = 12 else
"000000000000" when X = 176 AND Y = 12 else
"000000000000" when X = 177 AND Y = 12 else
"000000000000" when X = 178 AND Y = 12 else
"000000000000" when X = 179 AND Y = 12 else
"000000000000" when X = 180 AND Y = 12 else
"000000000000" when X = 181 AND Y = 12 else
"000000000000" when X = 182 AND Y = 12 else
"000000000000" when X = 183 AND Y = 12 else
"000000000000" when X = 184 AND Y = 12 else
"000000000000" when X = 185 AND Y = 12 else
"000000000000" when X = 186 AND Y = 12 else
"000000000000" when X = 187 AND Y = 12 else
"000000000000" when X = 188 AND Y = 12 else
"000000000000" when X = 189 AND Y = 12 else
"000000000000" when X = 190 AND Y = 12 else
"000000000000" when X = 191 AND Y = 12 else
"000000000000" when X = 192 AND Y = 12 else
"000000000000" when X = 193 AND Y = 12 else
"000000000000" when X = 194 AND Y = 12 else
"000000000000" when X = 195 AND Y = 12 else
"000000000000" when X = 196 AND Y = 12 else
"000000000000" when X = 197 AND Y = 12 else
"000000000000" when X = 198 AND Y = 12 else
"000000000000" when X = 199 AND Y = 12 else
"000000000000" when X = 200 AND Y = 12 else
"000000000000" when X = 201 AND Y = 12 else
"000000000000" when X = 202 AND Y = 12 else
"000000000000" when X = 203 AND Y = 12 else
"000000000000" when X = 204 AND Y = 12 else
"000000000000" when X = 205 AND Y = 12 else
"000000000000" when X = 206 AND Y = 12 else
"000000000000" when X = 207 AND Y = 12 else
"000000000000" when X = 208 AND Y = 12 else
"000000000000" when X = 209 AND Y = 12 else
"000000000000" when X = 210 AND Y = 12 else
"000000000000" when X = 211 AND Y = 12 else
"000000000000" when X = 212 AND Y = 12 else
"000000000000" when X = 213 AND Y = 12 else
"000000000000" when X = 214 AND Y = 12 else
"000000000000" when X = 215 AND Y = 12 else
"000000000000" when X = 216 AND Y = 12 else
"000000000000" when X = 217 AND Y = 12 else
"000000000000" when X = 218 AND Y = 12 else
"000000000000" when X = 219 AND Y = 12 else
"000000000000" when X = 220 AND Y = 12 else
"000000000000" when X = 221 AND Y = 12 else
"000000000000" when X = 222 AND Y = 12 else
"000000000000" when X = 223 AND Y = 12 else
"000000000000" when X = 224 AND Y = 12 else
"000000000000" when X = 225 AND Y = 12 else
"000000000000" when X = 226 AND Y = 12 else
"000000000000" when X = 227 AND Y = 12 else
"000000000000" when X = 228 AND Y = 12 else
"000000000000" when X = 229 AND Y = 12 else
"000000000000" when X = 230 AND Y = 12 else
"000000000000" when X = 231 AND Y = 12 else
"000000000000" when X = 232 AND Y = 12 else
"000000000000" when X = 233 AND Y = 12 else
"000000000000" when X = 234 AND Y = 12 else
"000000000000" when X = 235 AND Y = 12 else
"000000000000" when X = 236 AND Y = 12 else
"000000000000" when X = 237 AND Y = 12 else
"000000000000" when X = 238 AND Y = 12 else
"000000000000" when X = 239 AND Y = 12 else
"000000000000" when X = 240 AND Y = 12 else
"000000000000" when X = 241 AND Y = 12 else
"000000000000" when X = 242 AND Y = 12 else
"000000000000" when X = 243 AND Y = 12 else
"000000000000" when X = 244 AND Y = 12 else
"000000000000" when X = 245 AND Y = 12 else
"000000000000" when X = 246 AND Y = 12 else
"000000000000" when X = 247 AND Y = 12 else
"000000000000" when X = 248 AND Y = 12 else
"000000000000" when X = 249 AND Y = 12 else
"000000000000" when X = 250 AND Y = 12 else
"000000000000" when X = 251 AND Y = 12 else
"000000000000" when X = 252 AND Y = 12 else
"000000000000" when X = 253 AND Y = 12 else
"000000000000" when X = 254 AND Y = 12 else
"000000000000" when X = 255 AND Y = 12 else
"000000000000" when X = 256 AND Y = 12 else
"000000000000" when X = 257 AND Y = 12 else
"000000000000" when X = 258 AND Y = 12 else
"000000000000" when X = 259 AND Y = 12 else
"000000000000" when X = 260 AND Y = 12 else
"000000000000" when X = 261 AND Y = 12 else
"000000000000" when X = 262 AND Y = 12 else
"000000000000" when X = 263 AND Y = 12 else
"000000000000" when X = 264 AND Y = 12 else
"000000000000" when X = 265 AND Y = 12 else
"000000000000" when X = 266 AND Y = 12 else
"000000000000" when X = 267 AND Y = 12 else
"000000000000" when X = 268 AND Y = 12 else
"000000000000" when X = 269 AND Y = 12 else
"000000000000" when X = 270 AND Y = 12 else
"000000000000" when X = 271 AND Y = 12 else
"000000000000" when X = 272 AND Y = 12 else
"000000000000" when X = 273 AND Y = 12 else
"000000000000" when X = 274 AND Y = 12 else
"000000000000" when X = 275 AND Y = 12 else
"000000000000" when X = 276 AND Y = 12 else
"000000000000" when X = 277 AND Y = 12 else
"000000000000" when X = 278 AND Y = 12 else
"000000000000" when X = 279 AND Y = 12 else
"000000000000" when X = 280 AND Y = 12 else
"000000000000" when X = 281 AND Y = 12 else
"000000000000" when X = 282 AND Y = 12 else
"000000000000" when X = 283 AND Y = 12 else
"000000000000" when X = 284 AND Y = 12 else
"000000000000" when X = 285 AND Y = 12 else
"000000000000" when X = 286 AND Y = 12 else
"000000000000" when X = 287 AND Y = 12 else
"000000000000" when X = 288 AND Y = 12 else
"000000000000" when X = 289 AND Y = 12 else
"000000000000" when X = 290 AND Y = 12 else
"000000000000" when X = 291 AND Y = 12 else
"000000000000" when X = 292 AND Y = 12 else
"000000000000" when X = 293 AND Y = 12 else
"000000000000" when X = 294 AND Y = 12 else
"000000000000" when X = 295 AND Y = 12 else
"000000000000" when X = 296 AND Y = 12 else
"000000000000" when X = 297 AND Y = 12 else
"000000000000" when X = 298 AND Y = 12 else
"000000000000" when X = 299 AND Y = 12 else
"000000000000" when X = 300 AND Y = 12 else
"000000000000" when X = 301 AND Y = 12 else
"000000000000" when X = 302 AND Y = 12 else
"000000000000" when X = 303 AND Y = 12 else
"000000000000" when X = 304 AND Y = 12 else
"000000000000" when X = 305 AND Y = 12 else
"000000000000" when X = 306 AND Y = 12 else
"000000000000" when X = 307 AND Y = 12 else
"000000000000" when X = 308 AND Y = 12 else
"000000000000" when X = 309 AND Y = 12 else
"000000000000" when X = 310 AND Y = 12 else
"000000000000" when X = 311 AND Y = 12 else
"000000000000" when X = 312 AND Y = 12 else
"000000000000" when X = 313 AND Y = 12 else
"000000000000" when X = 314 AND Y = 12 else
"000000000000" when X = 315 AND Y = 12 else
"000000000000" when X = 316 AND Y = 12 else
"000000000000" when X = 317 AND Y = 12 else
"000000000000" when X = 318 AND Y = 12 else
"000000000000" when X = 319 AND Y = 12 else
"000000000000" when X = 320 AND Y = 12 else
"000000000000" when X = 321 AND Y = 12 else
"000000000000" when X = 322 AND Y = 12 else
"000000000000" when X = 323 AND Y = 12 else
"000000000000" when X = 324 AND Y = 12 else
"000000000000" when X = 0 AND Y = 13 else
"000000000000" when X = 1 AND Y = 13 else
"000000000000" when X = 2 AND Y = 13 else
"000000000000" when X = 3 AND Y = 13 else
"000000000000" when X = 4 AND Y = 13 else
"000000000000" when X = 5 AND Y = 13 else
"000000000000" when X = 6 AND Y = 13 else
"000000000000" when X = 7 AND Y = 13 else
"000000000000" when X = 8 AND Y = 13 else
"000000000000" when X = 9 AND Y = 13 else
"000000000000" when X = 10 AND Y = 13 else
"000000000000" when X = 11 AND Y = 13 else
"000000000000" when X = 12 AND Y = 13 else
"000000000000" when X = 13 AND Y = 13 else
"000000000000" when X = 14 AND Y = 13 else
"000000000000" when X = 15 AND Y = 13 else
"000000000000" when X = 16 AND Y = 13 else
"000000000000" when X = 17 AND Y = 13 else
"000000000000" when X = 18 AND Y = 13 else
"000000000000" when X = 19 AND Y = 13 else
"000000000000" when X = 20 AND Y = 13 else
"000000000000" when X = 21 AND Y = 13 else
"000000000000" when X = 22 AND Y = 13 else
"000000000000" when X = 23 AND Y = 13 else
"000000000000" when X = 24 AND Y = 13 else
"000000000000" when X = 25 AND Y = 13 else
"000000000000" when X = 26 AND Y = 13 else
"000000000000" when X = 27 AND Y = 13 else
"000000000000" when X = 28 AND Y = 13 else
"000000000000" when X = 29 AND Y = 13 else
"000000000000" when X = 30 AND Y = 13 else
"000000000000" when X = 31 AND Y = 13 else
"000000000000" when X = 32 AND Y = 13 else
"000000000000" when X = 33 AND Y = 13 else
"000000000000" when X = 34 AND Y = 13 else
"000000000000" when X = 35 AND Y = 13 else
"000000000000" when X = 36 AND Y = 13 else
"000000000000" when X = 37 AND Y = 13 else
"000000000000" when X = 38 AND Y = 13 else
"000000000000" when X = 39 AND Y = 13 else
"100010011101" when X = 40 AND Y = 13 else
"100010011101" when X = 41 AND Y = 13 else
"100010011101" when X = 42 AND Y = 13 else
"100010011101" when X = 43 AND Y = 13 else
"100010011101" when X = 44 AND Y = 13 else
"100010011101" when X = 45 AND Y = 13 else
"100010011101" when X = 46 AND Y = 13 else
"100010011101" when X = 47 AND Y = 13 else
"100010011101" when X = 48 AND Y = 13 else
"100010011101" when X = 49 AND Y = 13 else
"110111011111" when X = 50 AND Y = 13 else
"110111011111" when X = 51 AND Y = 13 else
"110111011111" when X = 52 AND Y = 13 else
"110111011111" when X = 53 AND Y = 13 else
"110111011111" when X = 54 AND Y = 13 else
"110111011111" when X = 55 AND Y = 13 else
"110111011111" when X = 56 AND Y = 13 else
"110111011111" when X = 57 AND Y = 13 else
"110111011111" when X = 58 AND Y = 13 else
"110111011111" when X = 59 AND Y = 13 else
"110111011111" when X = 60 AND Y = 13 else
"110111011111" when X = 61 AND Y = 13 else
"110111011111" when X = 62 AND Y = 13 else
"110111011111" when X = 63 AND Y = 13 else
"110111011111" when X = 64 AND Y = 13 else
"110111011111" when X = 65 AND Y = 13 else
"110111011111" when X = 66 AND Y = 13 else
"110111011111" when X = 67 AND Y = 13 else
"110111011111" when X = 68 AND Y = 13 else
"110111011111" when X = 69 AND Y = 13 else
"111111111111" when X = 70 AND Y = 13 else
"111111111111" when X = 71 AND Y = 13 else
"111111111111" when X = 72 AND Y = 13 else
"111111111111" when X = 73 AND Y = 13 else
"111111111111" when X = 74 AND Y = 13 else
"111111111111" when X = 75 AND Y = 13 else
"111111111111" when X = 76 AND Y = 13 else
"111111111111" when X = 77 AND Y = 13 else
"111111111111" when X = 78 AND Y = 13 else
"111111111111" when X = 79 AND Y = 13 else
"111111111111" when X = 80 AND Y = 13 else
"111111111111" when X = 81 AND Y = 13 else
"111111111111" when X = 82 AND Y = 13 else
"111111111111" when X = 83 AND Y = 13 else
"111111111111" when X = 84 AND Y = 13 else
"111111111111" when X = 85 AND Y = 13 else
"111111111111" when X = 86 AND Y = 13 else
"111111111111" when X = 87 AND Y = 13 else
"111111111111" when X = 88 AND Y = 13 else
"111111111111" when X = 89 AND Y = 13 else
"111111111111" when X = 90 AND Y = 13 else
"111111111111" when X = 91 AND Y = 13 else
"111111111111" when X = 92 AND Y = 13 else
"111111111111" when X = 93 AND Y = 13 else
"111111111111" when X = 94 AND Y = 13 else
"111111111111" when X = 95 AND Y = 13 else
"111111111111" when X = 96 AND Y = 13 else
"111111111111" when X = 97 AND Y = 13 else
"111111111111" when X = 98 AND Y = 13 else
"111111111111" when X = 99 AND Y = 13 else
"111111111111" when X = 100 AND Y = 13 else
"111111111111" when X = 101 AND Y = 13 else
"111111111111" when X = 102 AND Y = 13 else
"111111111111" when X = 103 AND Y = 13 else
"111111111111" when X = 104 AND Y = 13 else
"111111111111" when X = 105 AND Y = 13 else
"111111111111" when X = 106 AND Y = 13 else
"111111111111" when X = 107 AND Y = 13 else
"111111111111" when X = 108 AND Y = 13 else
"111111111111" when X = 109 AND Y = 13 else
"111111111111" when X = 110 AND Y = 13 else
"111111111111" when X = 111 AND Y = 13 else
"111111111111" when X = 112 AND Y = 13 else
"111111111111" when X = 113 AND Y = 13 else
"111111111111" when X = 114 AND Y = 13 else
"111111111111" when X = 115 AND Y = 13 else
"111111111111" when X = 116 AND Y = 13 else
"111111111111" when X = 117 AND Y = 13 else
"111111111111" when X = 118 AND Y = 13 else
"111111111111" when X = 119 AND Y = 13 else
"111111111111" when X = 120 AND Y = 13 else
"111111111111" when X = 121 AND Y = 13 else
"111111111111" when X = 122 AND Y = 13 else
"111111111111" when X = 123 AND Y = 13 else
"111111111111" when X = 124 AND Y = 13 else
"111111111111" when X = 125 AND Y = 13 else
"111111111111" when X = 126 AND Y = 13 else
"111111111111" when X = 127 AND Y = 13 else
"111111111111" when X = 128 AND Y = 13 else
"111111111111" when X = 129 AND Y = 13 else
"111111111111" when X = 130 AND Y = 13 else
"111111111111" when X = 131 AND Y = 13 else
"111111111111" when X = 132 AND Y = 13 else
"111111111111" when X = 133 AND Y = 13 else
"111111111111" when X = 134 AND Y = 13 else
"111111111111" when X = 135 AND Y = 13 else
"111111111111" when X = 136 AND Y = 13 else
"111111111111" when X = 137 AND Y = 13 else
"111111111111" when X = 138 AND Y = 13 else
"111111111111" when X = 139 AND Y = 13 else
"111111111111" when X = 140 AND Y = 13 else
"111111111111" when X = 141 AND Y = 13 else
"111111111111" when X = 142 AND Y = 13 else
"111111111111" when X = 143 AND Y = 13 else
"111111111111" when X = 144 AND Y = 13 else
"111111111111" when X = 145 AND Y = 13 else
"111111111111" when X = 146 AND Y = 13 else
"111111111111" when X = 147 AND Y = 13 else
"111111111111" when X = 148 AND Y = 13 else
"111111111111" when X = 149 AND Y = 13 else
"000000000000" when X = 150 AND Y = 13 else
"000000000000" when X = 151 AND Y = 13 else
"000000000000" when X = 152 AND Y = 13 else
"000000000000" when X = 153 AND Y = 13 else
"000000000000" when X = 154 AND Y = 13 else
"000000000000" when X = 155 AND Y = 13 else
"000000000000" when X = 156 AND Y = 13 else
"000000000000" when X = 157 AND Y = 13 else
"000000000000" when X = 158 AND Y = 13 else
"000000000000" when X = 159 AND Y = 13 else
"000000000000" when X = 160 AND Y = 13 else
"000000000000" when X = 161 AND Y = 13 else
"000000000000" when X = 162 AND Y = 13 else
"000000000000" when X = 163 AND Y = 13 else
"000000000000" when X = 164 AND Y = 13 else
"000000000000" when X = 165 AND Y = 13 else
"000000000000" when X = 166 AND Y = 13 else
"000000000000" when X = 167 AND Y = 13 else
"000000000000" when X = 168 AND Y = 13 else
"000000000000" when X = 169 AND Y = 13 else
"000000000000" when X = 170 AND Y = 13 else
"000000000000" when X = 171 AND Y = 13 else
"000000000000" when X = 172 AND Y = 13 else
"000000000000" when X = 173 AND Y = 13 else
"000000000000" when X = 174 AND Y = 13 else
"000000000000" when X = 175 AND Y = 13 else
"000000000000" when X = 176 AND Y = 13 else
"000000000000" when X = 177 AND Y = 13 else
"000000000000" when X = 178 AND Y = 13 else
"000000000000" when X = 179 AND Y = 13 else
"000000000000" when X = 180 AND Y = 13 else
"000000000000" when X = 181 AND Y = 13 else
"000000000000" when X = 182 AND Y = 13 else
"000000000000" when X = 183 AND Y = 13 else
"000000000000" when X = 184 AND Y = 13 else
"000000000000" when X = 185 AND Y = 13 else
"000000000000" when X = 186 AND Y = 13 else
"000000000000" when X = 187 AND Y = 13 else
"000000000000" when X = 188 AND Y = 13 else
"000000000000" when X = 189 AND Y = 13 else
"000000000000" when X = 190 AND Y = 13 else
"000000000000" when X = 191 AND Y = 13 else
"000000000000" when X = 192 AND Y = 13 else
"000000000000" when X = 193 AND Y = 13 else
"000000000000" when X = 194 AND Y = 13 else
"000000000000" when X = 195 AND Y = 13 else
"000000000000" when X = 196 AND Y = 13 else
"000000000000" when X = 197 AND Y = 13 else
"000000000000" when X = 198 AND Y = 13 else
"000000000000" when X = 199 AND Y = 13 else
"000000000000" when X = 200 AND Y = 13 else
"000000000000" when X = 201 AND Y = 13 else
"000000000000" when X = 202 AND Y = 13 else
"000000000000" when X = 203 AND Y = 13 else
"000000000000" when X = 204 AND Y = 13 else
"000000000000" when X = 205 AND Y = 13 else
"000000000000" when X = 206 AND Y = 13 else
"000000000000" when X = 207 AND Y = 13 else
"000000000000" when X = 208 AND Y = 13 else
"000000000000" when X = 209 AND Y = 13 else
"000000000000" when X = 210 AND Y = 13 else
"000000000000" when X = 211 AND Y = 13 else
"000000000000" when X = 212 AND Y = 13 else
"000000000000" when X = 213 AND Y = 13 else
"000000000000" when X = 214 AND Y = 13 else
"000000000000" when X = 215 AND Y = 13 else
"000000000000" when X = 216 AND Y = 13 else
"000000000000" when X = 217 AND Y = 13 else
"000000000000" when X = 218 AND Y = 13 else
"000000000000" when X = 219 AND Y = 13 else
"000000000000" when X = 220 AND Y = 13 else
"000000000000" when X = 221 AND Y = 13 else
"000000000000" when X = 222 AND Y = 13 else
"000000000000" when X = 223 AND Y = 13 else
"000000000000" when X = 224 AND Y = 13 else
"000000000000" when X = 225 AND Y = 13 else
"000000000000" when X = 226 AND Y = 13 else
"000000000000" when X = 227 AND Y = 13 else
"000000000000" when X = 228 AND Y = 13 else
"000000000000" when X = 229 AND Y = 13 else
"000000000000" when X = 230 AND Y = 13 else
"000000000000" when X = 231 AND Y = 13 else
"000000000000" when X = 232 AND Y = 13 else
"000000000000" when X = 233 AND Y = 13 else
"000000000000" when X = 234 AND Y = 13 else
"000000000000" when X = 235 AND Y = 13 else
"000000000000" when X = 236 AND Y = 13 else
"000000000000" when X = 237 AND Y = 13 else
"000000000000" when X = 238 AND Y = 13 else
"000000000000" when X = 239 AND Y = 13 else
"000000000000" when X = 240 AND Y = 13 else
"000000000000" when X = 241 AND Y = 13 else
"000000000000" when X = 242 AND Y = 13 else
"000000000000" when X = 243 AND Y = 13 else
"000000000000" when X = 244 AND Y = 13 else
"000000000000" when X = 245 AND Y = 13 else
"000000000000" when X = 246 AND Y = 13 else
"000000000000" when X = 247 AND Y = 13 else
"000000000000" when X = 248 AND Y = 13 else
"000000000000" when X = 249 AND Y = 13 else
"000000000000" when X = 250 AND Y = 13 else
"000000000000" when X = 251 AND Y = 13 else
"000000000000" when X = 252 AND Y = 13 else
"000000000000" when X = 253 AND Y = 13 else
"000000000000" when X = 254 AND Y = 13 else
"000000000000" when X = 255 AND Y = 13 else
"000000000000" when X = 256 AND Y = 13 else
"000000000000" when X = 257 AND Y = 13 else
"000000000000" when X = 258 AND Y = 13 else
"000000000000" when X = 259 AND Y = 13 else
"000000000000" when X = 260 AND Y = 13 else
"000000000000" when X = 261 AND Y = 13 else
"000000000000" when X = 262 AND Y = 13 else
"000000000000" when X = 263 AND Y = 13 else
"000000000000" when X = 264 AND Y = 13 else
"000000000000" when X = 265 AND Y = 13 else
"000000000000" when X = 266 AND Y = 13 else
"000000000000" when X = 267 AND Y = 13 else
"000000000000" when X = 268 AND Y = 13 else
"000000000000" when X = 269 AND Y = 13 else
"000000000000" when X = 270 AND Y = 13 else
"000000000000" when X = 271 AND Y = 13 else
"000000000000" when X = 272 AND Y = 13 else
"000000000000" when X = 273 AND Y = 13 else
"000000000000" when X = 274 AND Y = 13 else
"000000000000" when X = 275 AND Y = 13 else
"000000000000" when X = 276 AND Y = 13 else
"000000000000" when X = 277 AND Y = 13 else
"000000000000" when X = 278 AND Y = 13 else
"000000000000" when X = 279 AND Y = 13 else
"000000000000" when X = 280 AND Y = 13 else
"000000000000" when X = 281 AND Y = 13 else
"000000000000" when X = 282 AND Y = 13 else
"000000000000" when X = 283 AND Y = 13 else
"000000000000" when X = 284 AND Y = 13 else
"000000000000" when X = 285 AND Y = 13 else
"000000000000" when X = 286 AND Y = 13 else
"000000000000" when X = 287 AND Y = 13 else
"000000000000" when X = 288 AND Y = 13 else
"000000000000" when X = 289 AND Y = 13 else
"000000000000" when X = 290 AND Y = 13 else
"000000000000" when X = 291 AND Y = 13 else
"000000000000" when X = 292 AND Y = 13 else
"000000000000" when X = 293 AND Y = 13 else
"000000000000" when X = 294 AND Y = 13 else
"000000000000" when X = 295 AND Y = 13 else
"000000000000" when X = 296 AND Y = 13 else
"000000000000" when X = 297 AND Y = 13 else
"000000000000" when X = 298 AND Y = 13 else
"000000000000" when X = 299 AND Y = 13 else
"000000000000" when X = 300 AND Y = 13 else
"000000000000" when X = 301 AND Y = 13 else
"000000000000" when X = 302 AND Y = 13 else
"000000000000" when X = 303 AND Y = 13 else
"000000000000" when X = 304 AND Y = 13 else
"000000000000" when X = 305 AND Y = 13 else
"000000000000" when X = 306 AND Y = 13 else
"000000000000" when X = 307 AND Y = 13 else
"000000000000" when X = 308 AND Y = 13 else
"000000000000" when X = 309 AND Y = 13 else
"000000000000" when X = 310 AND Y = 13 else
"000000000000" when X = 311 AND Y = 13 else
"000000000000" when X = 312 AND Y = 13 else
"000000000000" when X = 313 AND Y = 13 else
"000000000000" when X = 314 AND Y = 13 else
"000000000000" when X = 315 AND Y = 13 else
"000000000000" when X = 316 AND Y = 13 else
"000000000000" when X = 317 AND Y = 13 else
"000000000000" when X = 318 AND Y = 13 else
"000000000000" when X = 319 AND Y = 13 else
"000000000000" when X = 320 AND Y = 13 else
"000000000000" when X = 321 AND Y = 13 else
"000000000000" when X = 322 AND Y = 13 else
"000000000000" when X = 323 AND Y = 13 else
"000000000000" when X = 324 AND Y = 13 else
"000000000000" when X = 0 AND Y = 14 else
"000000000000" when X = 1 AND Y = 14 else
"000000000000" when X = 2 AND Y = 14 else
"000000000000" when X = 3 AND Y = 14 else
"000000000000" when X = 4 AND Y = 14 else
"000000000000" when X = 5 AND Y = 14 else
"000000000000" when X = 6 AND Y = 14 else
"000000000000" when X = 7 AND Y = 14 else
"000000000000" when X = 8 AND Y = 14 else
"000000000000" when X = 9 AND Y = 14 else
"000000000000" when X = 10 AND Y = 14 else
"000000000000" when X = 11 AND Y = 14 else
"000000000000" when X = 12 AND Y = 14 else
"000000000000" when X = 13 AND Y = 14 else
"000000000000" when X = 14 AND Y = 14 else
"000000000000" when X = 15 AND Y = 14 else
"000000000000" when X = 16 AND Y = 14 else
"000000000000" when X = 17 AND Y = 14 else
"000000000000" when X = 18 AND Y = 14 else
"000000000000" when X = 19 AND Y = 14 else
"000000000000" when X = 20 AND Y = 14 else
"000000000000" when X = 21 AND Y = 14 else
"000000000000" when X = 22 AND Y = 14 else
"000000000000" when X = 23 AND Y = 14 else
"000000000000" when X = 24 AND Y = 14 else
"000000000000" when X = 25 AND Y = 14 else
"000000000000" when X = 26 AND Y = 14 else
"000000000000" when X = 27 AND Y = 14 else
"000000000000" when X = 28 AND Y = 14 else
"000000000000" when X = 29 AND Y = 14 else
"000000000000" when X = 30 AND Y = 14 else
"000000000000" when X = 31 AND Y = 14 else
"000000000000" when X = 32 AND Y = 14 else
"000000000000" when X = 33 AND Y = 14 else
"000000000000" when X = 34 AND Y = 14 else
"000000000000" when X = 35 AND Y = 14 else
"000000000000" when X = 36 AND Y = 14 else
"000000000000" when X = 37 AND Y = 14 else
"000000000000" when X = 38 AND Y = 14 else
"000000000000" when X = 39 AND Y = 14 else
"100010011101" when X = 40 AND Y = 14 else
"100010011101" when X = 41 AND Y = 14 else
"100010011101" when X = 42 AND Y = 14 else
"100010011101" when X = 43 AND Y = 14 else
"100010011101" when X = 44 AND Y = 14 else
"100010011101" when X = 45 AND Y = 14 else
"100010011101" when X = 46 AND Y = 14 else
"100010011101" when X = 47 AND Y = 14 else
"100010011101" when X = 48 AND Y = 14 else
"100010011101" when X = 49 AND Y = 14 else
"110111011111" when X = 50 AND Y = 14 else
"110111011111" when X = 51 AND Y = 14 else
"110111011111" when X = 52 AND Y = 14 else
"110111011111" when X = 53 AND Y = 14 else
"110111011111" when X = 54 AND Y = 14 else
"110111011111" when X = 55 AND Y = 14 else
"110111011111" when X = 56 AND Y = 14 else
"110111011111" when X = 57 AND Y = 14 else
"110111011111" when X = 58 AND Y = 14 else
"110111011111" when X = 59 AND Y = 14 else
"110111011111" when X = 60 AND Y = 14 else
"110111011111" when X = 61 AND Y = 14 else
"110111011111" when X = 62 AND Y = 14 else
"110111011111" when X = 63 AND Y = 14 else
"110111011111" when X = 64 AND Y = 14 else
"110111011111" when X = 65 AND Y = 14 else
"110111011111" when X = 66 AND Y = 14 else
"110111011111" when X = 67 AND Y = 14 else
"110111011111" when X = 68 AND Y = 14 else
"110111011111" when X = 69 AND Y = 14 else
"111111111111" when X = 70 AND Y = 14 else
"111111111111" when X = 71 AND Y = 14 else
"111111111111" when X = 72 AND Y = 14 else
"111111111111" when X = 73 AND Y = 14 else
"111111111111" when X = 74 AND Y = 14 else
"111111111111" when X = 75 AND Y = 14 else
"111111111111" when X = 76 AND Y = 14 else
"111111111111" when X = 77 AND Y = 14 else
"111111111111" when X = 78 AND Y = 14 else
"111111111111" when X = 79 AND Y = 14 else
"111111111111" when X = 80 AND Y = 14 else
"111111111111" when X = 81 AND Y = 14 else
"111111111111" when X = 82 AND Y = 14 else
"111111111111" when X = 83 AND Y = 14 else
"111111111111" when X = 84 AND Y = 14 else
"111111111111" when X = 85 AND Y = 14 else
"111111111111" when X = 86 AND Y = 14 else
"111111111111" when X = 87 AND Y = 14 else
"111111111111" when X = 88 AND Y = 14 else
"111111111111" when X = 89 AND Y = 14 else
"111111111111" when X = 90 AND Y = 14 else
"111111111111" when X = 91 AND Y = 14 else
"111111111111" when X = 92 AND Y = 14 else
"111111111111" when X = 93 AND Y = 14 else
"111111111111" when X = 94 AND Y = 14 else
"111111111111" when X = 95 AND Y = 14 else
"111111111111" when X = 96 AND Y = 14 else
"111111111111" when X = 97 AND Y = 14 else
"111111111111" when X = 98 AND Y = 14 else
"111111111111" when X = 99 AND Y = 14 else
"111111111111" when X = 100 AND Y = 14 else
"111111111111" when X = 101 AND Y = 14 else
"111111111111" when X = 102 AND Y = 14 else
"111111111111" when X = 103 AND Y = 14 else
"111111111111" when X = 104 AND Y = 14 else
"111111111111" when X = 105 AND Y = 14 else
"111111111111" when X = 106 AND Y = 14 else
"111111111111" when X = 107 AND Y = 14 else
"111111111111" when X = 108 AND Y = 14 else
"111111111111" when X = 109 AND Y = 14 else
"111111111111" when X = 110 AND Y = 14 else
"111111111111" when X = 111 AND Y = 14 else
"111111111111" when X = 112 AND Y = 14 else
"111111111111" when X = 113 AND Y = 14 else
"111111111111" when X = 114 AND Y = 14 else
"111111111111" when X = 115 AND Y = 14 else
"111111111111" when X = 116 AND Y = 14 else
"111111111111" when X = 117 AND Y = 14 else
"111111111111" when X = 118 AND Y = 14 else
"111111111111" when X = 119 AND Y = 14 else
"111111111111" when X = 120 AND Y = 14 else
"111111111111" when X = 121 AND Y = 14 else
"111111111111" when X = 122 AND Y = 14 else
"111111111111" when X = 123 AND Y = 14 else
"111111111111" when X = 124 AND Y = 14 else
"111111111111" when X = 125 AND Y = 14 else
"111111111111" when X = 126 AND Y = 14 else
"111111111111" when X = 127 AND Y = 14 else
"111111111111" when X = 128 AND Y = 14 else
"111111111111" when X = 129 AND Y = 14 else
"111111111111" when X = 130 AND Y = 14 else
"111111111111" when X = 131 AND Y = 14 else
"111111111111" when X = 132 AND Y = 14 else
"111111111111" when X = 133 AND Y = 14 else
"111111111111" when X = 134 AND Y = 14 else
"111111111111" when X = 135 AND Y = 14 else
"111111111111" when X = 136 AND Y = 14 else
"111111111111" when X = 137 AND Y = 14 else
"111111111111" when X = 138 AND Y = 14 else
"111111111111" when X = 139 AND Y = 14 else
"111111111111" when X = 140 AND Y = 14 else
"111111111111" when X = 141 AND Y = 14 else
"111111111111" when X = 142 AND Y = 14 else
"111111111111" when X = 143 AND Y = 14 else
"111111111111" when X = 144 AND Y = 14 else
"111111111111" when X = 145 AND Y = 14 else
"111111111111" when X = 146 AND Y = 14 else
"111111111111" when X = 147 AND Y = 14 else
"111111111111" when X = 148 AND Y = 14 else
"111111111111" when X = 149 AND Y = 14 else
"000000000000" when X = 150 AND Y = 14 else
"000000000000" when X = 151 AND Y = 14 else
"000000000000" when X = 152 AND Y = 14 else
"000000000000" when X = 153 AND Y = 14 else
"000000000000" when X = 154 AND Y = 14 else
"000000000000" when X = 155 AND Y = 14 else
"000000000000" when X = 156 AND Y = 14 else
"000000000000" when X = 157 AND Y = 14 else
"000000000000" when X = 158 AND Y = 14 else
"000000000000" when X = 159 AND Y = 14 else
"000000000000" when X = 160 AND Y = 14 else
"000000000000" when X = 161 AND Y = 14 else
"000000000000" when X = 162 AND Y = 14 else
"000000000000" when X = 163 AND Y = 14 else
"000000000000" when X = 164 AND Y = 14 else
"000000000000" when X = 165 AND Y = 14 else
"000000000000" when X = 166 AND Y = 14 else
"000000000000" when X = 167 AND Y = 14 else
"000000000000" when X = 168 AND Y = 14 else
"000000000000" when X = 169 AND Y = 14 else
"000000000000" when X = 170 AND Y = 14 else
"000000000000" when X = 171 AND Y = 14 else
"000000000000" when X = 172 AND Y = 14 else
"000000000000" when X = 173 AND Y = 14 else
"000000000000" when X = 174 AND Y = 14 else
"000000000000" when X = 175 AND Y = 14 else
"000000000000" when X = 176 AND Y = 14 else
"000000000000" when X = 177 AND Y = 14 else
"000000000000" when X = 178 AND Y = 14 else
"000000000000" when X = 179 AND Y = 14 else
"000000000000" when X = 180 AND Y = 14 else
"000000000000" when X = 181 AND Y = 14 else
"000000000000" when X = 182 AND Y = 14 else
"000000000000" when X = 183 AND Y = 14 else
"000000000000" when X = 184 AND Y = 14 else
"000000000000" when X = 185 AND Y = 14 else
"000000000000" when X = 186 AND Y = 14 else
"000000000000" when X = 187 AND Y = 14 else
"000000000000" when X = 188 AND Y = 14 else
"000000000000" when X = 189 AND Y = 14 else
"000000000000" when X = 190 AND Y = 14 else
"000000000000" when X = 191 AND Y = 14 else
"000000000000" when X = 192 AND Y = 14 else
"000000000000" when X = 193 AND Y = 14 else
"000000000000" when X = 194 AND Y = 14 else
"000000000000" when X = 195 AND Y = 14 else
"000000000000" when X = 196 AND Y = 14 else
"000000000000" when X = 197 AND Y = 14 else
"000000000000" when X = 198 AND Y = 14 else
"000000000000" when X = 199 AND Y = 14 else
"000000000000" when X = 200 AND Y = 14 else
"000000000000" when X = 201 AND Y = 14 else
"000000000000" when X = 202 AND Y = 14 else
"000000000000" when X = 203 AND Y = 14 else
"000000000000" when X = 204 AND Y = 14 else
"000000000000" when X = 205 AND Y = 14 else
"000000000000" when X = 206 AND Y = 14 else
"000000000000" when X = 207 AND Y = 14 else
"000000000000" when X = 208 AND Y = 14 else
"000000000000" when X = 209 AND Y = 14 else
"000000000000" when X = 210 AND Y = 14 else
"000000000000" when X = 211 AND Y = 14 else
"000000000000" when X = 212 AND Y = 14 else
"000000000000" when X = 213 AND Y = 14 else
"000000000000" when X = 214 AND Y = 14 else
"000000000000" when X = 215 AND Y = 14 else
"000000000000" when X = 216 AND Y = 14 else
"000000000000" when X = 217 AND Y = 14 else
"000000000000" when X = 218 AND Y = 14 else
"000000000000" when X = 219 AND Y = 14 else
"000000000000" when X = 220 AND Y = 14 else
"000000000000" when X = 221 AND Y = 14 else
"000000000000" when X = 222 AND Y = 14 else
"000000000000" when X = 223 AND Y = 14 else
"000000000000" when X = 224 AND Y = 14 else
"000000000000" when X = 225 AND Y = 14 else
"000000000000" when X = 226 AND Y = 14 else
"000000000000" when X = 227 AND Y = 14 else
"000000000000" when X = 228 AND Y = 14 else
"000000000000" when X = 229 AND Y = 14 else
"000000000000" when X = 230 AND Y = 14 else
"000000000000" when X = 231 AND Y = 14 else
"000000000000" when X = 232 AND Y = 14 else
"000000000000" when X = 233 AND Y = 14 else
"000000000000" when X = 234 AND Y = 14 else
"000000000000" when X = 235 AND Y = 14 else
"000000000000" when X = 236 AND Y = 14 else
"000000000000" when X = 237 AND Y = 14 else
"000000000000" when X = 238 AND Y = 14 else
"000000000000" when X = 239 AND Y = 14 else
"000000000000" when X = 240 AND Y = 14 else
"000000000000" when X = 241 AND Y = 14 else
"000000000000" when X = 242 AND Y = 14 else
"000000000000" when X = 243 AND Y = 14 else
"000000000000" when X = 244 AND Y = 14 else
"000000000000" when X = 245 AND Y = 14 else
"000000000000" when X = 246 AND Y = 14 else
"000000000000" when X = 247 AND Y = 14 else
"000000000000" when X = 248 AND Y = 14 else
"000000000000" when X = 249 AND Y = 14 else
"000000000000" when X = 250 AND Y = 14 else
"000000000000" when X = 251 AND Y = 14 else
"000000000000" when X = 252 AND Y = 14 else
"000000000000" when X = 253 AND Y = 14 else
"000000000000" when X = 254 AND Y = 14 else
"000000000000" when X = 255 AND Y = 14 else
"000000000000" when X = 256 AND Y = 14 else
"000000000000" when X = 257 AND Y = 14 else
"000000000000" when X = 258 AND Y = 14 else
"000000000000" when X = 259 AND Y = 14 else
"000000000000" when X = 260 AND Y = 14 else
"000000000000" when X = 261 AND Y = 14 else
"000000000000" when X = 262 AND Y = 14 else
"000000000000" when X = 263 AND Y = 14 else
"000000000000" when X = 264 AND Y = 14 else
"000000000000" when X = 265 AND Y = 14 else
"000000000000" when X = 266 AND Y = 14 else
"000000000000" when X = 267 AND Y = 14 else
"000000000000" when X = 268 AND Y = 14 else
"000000000000" when X = 269 AND Y = 14 else
"000000000000" when X = 270 AND Y = 14 else
"000000000000" when X = 271 AND Y = 14 else
"000000000000" when X = 272 AND Y = 14 else
"000000000000" when X = 273 AND Y = 14 else
"000000000000" when X = 274 AND Y = 14 else
"000000000000" when X = 275 AND Y = 14 else
"000000000000" when X = 276 AND Y = 14 else
"000000000000" when X = 277 AND Y = 14 else
"000000000000" when X = 278 AND Y = 14 else
"000000000000" when X = 279 AND Y = 14 else
"000000000000" when X = 280 AND Y = 14 else
"000000000000" when X = 281 AND Y = 14 else
"000000000000" when X = 282 AND Y = 14 else
"000000000000" when X = 283 AND Y = 14 else
"000000000000" when X = 284 AND Y = 14 else
"000000000000" when X = 285 AND Y = 14 else
"000000000000" when X = 286 AND Y = 14 else
"000000000000" when X = 287 AND Y = 14 else
"000000000000" when X = 288 AND Y = 14 else
"000000000000" when X = 289 AND Y = 14 else
"000000000000" when X = 290 AND Y = 14 else
"000000000000" when X = 291 AND Y = 14 else
"000000000000" when X = 292 AND Y = 14 else
"000000000000" when X = 293 AND Y = 14 else
"000000000000" when X = 294 AND Y = 14 else
"000000000000" when X = 295 AND Y = 14 else
"000000000000" when X = 296 AND Y = 14 else
"000000000000" when X = 297 AND Y = 14 else
"000000000000" when X = 298 AND Y = 14 else
"000000000000" when X = 299 AND Y = 14 else
"000000000000" when X = 300 AND Y = 14 else
"000000000000" when X = 301 AND Y = 14 else
"000000000000" when X = 302 AND Y = 14 else
"000000000000" when X = 303 AND Y = 14 else
"000000000000" when X = 304 AND Y = 14 else
"000000000000" when X = 305 AND Y = 14 else
"000000000000" when X = 306 AND Y = 14 else
"000000000000" when X = 307 AND Y = 14 else
"000000000000" when X = 308 AND Y = 14 else
"000000000000" when X = 309 AND Y = 14 else
"000000000000" when X = 310 AND Y = 14 else
"000000000000" when X = 311 AND Y = 14 else
"000000000000" when X = 312 AND Y = 14 else
"000000000000" when X = 313 AND Y = 14 else
"000000000000" when X = 314 AND Y = 14 else
"000000000000" when X = 315 AND Y = 14 else
"000000000000" when X = 316 AND Y = 14 else
"000000000000" when X = 317 AND Y = 14 else
"000000000000" when X = 318 AND Y = 14 else
"000000000000" when X = 319 AND Y = 14 else
"000000000000" when X = 320 AND Y = 14 else
"000000000000" when X = 321 AND Y = 14 else
"000000000000" when X = 322 AND Y = 14 else
"000000000000" when X = 323 AND Y = 14 else
"000000000000" when X = 324 AND Y = 14 else
"000000000000" when X = 0 AND Y = 15 else
"000000000000" when X = 1 AND Y = 15 else
"000000000000" when X = 2 AND Y = 15 else
"000000000000" when X = 3 AND Y = 15 else
"000000000000" when X = 4 AND Y = 15 else
"000000000000" when X = 5 AND Y = 15 else
"000000000000" when X = 6 AND Y = 15 else
"000000000000" when X = 7 AND Y = 15 else
"000000000000" when X = 8 AND Y = 15 else
"000000000000" when X = 9 AND Y = 15 else
"000000000000" when X = 10 AND Y = 15 else
"000000000000" when X = 11 AND Y = 15 else
"000000000000" when X = 12 AND Y = 15 else
"000000000000" when X = 13 AND Y = 15 else
"000000000000" when X = 14 AND Y = 15 else
"000000000000" when X = 15 AND Y = 15 else
"000000000000" when X = 16 AND Y = 15 else
"000000000000" when X = 17 AND Y = 15 else
"000000000000" when X = 18 AND Y = 15 else
"000000000000" when X = 19 AND Y = 15 else
"000000000000" when X = 20 AND Y = 15 else
"000000000000" when X = 21 AND Y = 15 else
"000000000000" when X = 22 AND Y = 15 else
"000000000000" when X = 23 AND Y = 15 else
"000000000000" when X = 24 AND Y = 15 else
"000000000000" when X = 25 AND Y = 15 else
"000000000000" when X = 26 AND Y = 15 else
"000000000000" when X = 27 AND Y = 15 else
"000000000000" when X = 28 AND Y = 15 else
"000000000000" when X = 29 AND Y = 15 else
"000000000000" when X = 30 AND Y = 15 else
"000000000000" when X = 31 AND Y = 15 else
"000000000000" when X = 32 AND Y = 15 else
"000000000000" when X = 33 AND Y = 15 else
"000000000000" when X = 34 AND Y = 15 else
"000000000000" when X = 35 AND Y = 15 else
"000000000000" when X = 36 AND Y = 15 else
"000000000000" when X = 37 AND Y = 15 else
"000000000000" when X = 38 AND Y = 15 else
"000000000000" when X = 39 AND Y = 15 else
"100010011101" when X = 40 AND Y = 15 else
"100010011101" when X = 41 AND Y = 15 else
"100010011101" when X = 42 AND Y = 15 else
"100010011101" when X = 43 AND Y = 15 else
"100010011101" when X = 44 AND Y = 15 else
"100010011101" when X = 45 AND Y = 15 else
"100010011101" when X = 46 AND Y = 15 else
"100010011101" when X = 47 AND Y = 15 else
"100010011101" when X = 48 AND Y = 15 else
"100010011101" when X = 49 AND Y = 15 else
"110111011111" when X = 50 AND Y = 15 else
"110111011111" when X = 51 AND Y = 15 else
"110111011111" when X = 52 AND Y = 15 else
"110111011111" when X = 53 AND Y = 15 else
"110111011111" when X = 54 AND Y = 15 else
"110111011111" when X = 55 AND Y = 15 else
"110111011111" when X = 56 AND Y = 15 else
"110111011111" when X = 57 AND Y = 15 else
"110111011111" when X = 58 AND Y = 15 else
"110111011111" when X = 59 AND Y = 15 else
"110111011111" when X = 60 AND Y = 15 else
"110111011111" when X = 61 AND Y = 15 else
"110111011111" when X = 62 AND Y = 15 else
"110111011111" when X = 63 AND Y = 15 else
"110111011111" when X = 64 AND Y = 15 else
"111111111111" when X = 65 AND Y = 15 else
"111111111111" when X = 66 AND Y = 15 else
"111111111111" when X = 67 AND Y = 15 else
"111111111111" when X = 68 AND Y = 15 else
"111111111111" when X = 69 AND Y = 15 else
"111111111111" when X = 70 AND Y = 15 else
"111111111111" when X = 71 AND Y = 15 else
"111111111111" when X = 72 AND Y = 15 else
"111111111111" when X = 73 AND Y = 15 else
"111111111111" when X = 74 AND Y = 15 else
"111111111111" when X = 75 AND Y = 15 else
"111111111111" when X = 76 AND Y = 15 else
"111111111111" when X = 77 AND Y = 15 else
"111111111111" when X = 78 AND Y = 15 else
"111111111111" when X = 79 AND Y = 15 else
"111111111111" when X = 80 AND Y = 15 else
"111111111111" when X = 81 AND Y = 15 else
"111111111111" when X = 82 AND Y = 15 else
"111111111111" when X = 83 AND Y = 15 else
"111111111111" when X = 84 AND Y = 15 else
"111111111111" when X = 85 AND Y = 15 else
"111111111111" when X = 86 AND Y = 15 else
"111111111111" when X = 87 AND Y = 15 else
"111111111111" when X = 88 AND Y = 15 else
"111111111111" when X = 89 AND Y = 15 else
"111111111111" when X = 90 AND Y = 15 else
"111111111111" when X = 91 AND Y = 15 else
"111111111111" when X = 92 AND Y = 15 else
"111111111111" when X = 93 AND Y = 15 else
"111111111111" when X = 94 AND Y = 15 else
"111111111111" when X = 95 AND Y = 15 else
"111111111111" when X = 96 AND Y = 15 else
"111111111111" when X = 97 AND Y = 15 else
"111111111111" when X = 98 AND Y = 15 else
"111111111111" when X = 99 AND Y = 15 else
"111111111111" when X = 100 AND Y = 15 else
"111111111111" when X = 101 AND Y = 15 else
"111111111111" when X = 102 AND Y = 15 else
"111111111111" when X = 103 AND Y = 15 else
"111111111111" when X = 104 AND Y = 15 else
"111111111111" when X = 105 AND Y = 15 else
"111111111111" when X = 106 AND Y = 15 else
"111111111111" when X = 107 AND Y = 15 else
"111111111111" when X = 108 AND Y = 15 else
"111111111111" when X = 109 AND Y = 15 else
"111111111111" when X = 110 AND Y = 15 else
"111111111111" when X = 111 AND Y = 15 else
"111111111111" when X = 112 AND Y = 15 else
"111111111111" when X = 113 AND Y = 15 else
"111111111111" when X = 114 AND Y = 15 else
"111111111111" when X = 115 AND Y = 15 else
"111111111111" when X = 116 AND Y = 15 else
"111111111111" when X = 117 AND Y = 15 else
"111111111111" when X = 118 AND Y = 15 else
"111111111111" when X = 119 AND Y = 15 else
"111111111111" when X = 120 AND Y = 15 else
"111111111111" when X = 121 AND Y = 15 else
"111111111111" when X = 122 AND Y = 15 else
"111111111111" when X = 123 AND Y = 15 else
"111111111111" when X = 124 AND Y = 15 else
"111111111111" when X = 125 AND Y = 15 else
"111111111111" when X = 126 AND Y = 15 else
"111111111111" when X = 127 AND Y = 15 else
"111111111111" when X = 128 AND Y = 15 else
"111111111111" when X = 129 AND Y = 15 else
"111111111111" when X = 130 AND Y = 15 else
"111111111111" when X = 131 AND Y = 15 else
"111111111111" when X = 132 AND Y = 15 else
"111111111111" when X = 133 AND Y = 15 else
"111111111111" when X = 134 AND Y = 15 else
"111111111111" when X = 135 AND Y = 15 else
"111111111111" when X = 136 AND Y = 15 else
"111111111111" when X = 137 AND Y = 15 else
"111111111111" when X = 138 AND Y = 15 else
"111111111111" when X = 139 AND Y = 15 else
"111111111111" when X = 140 AND Y = 15 else
"111111111111" when X = 141 AND Y = 15 else
"111111111111" when X = 142 AND Y = 15 else
"111111111111" when X = 143 AND Y = 15 else
"111111111111" when X = 144 AND Y = 15 else
"111111111111" when X = 145 AND Y = 15 else
"111111111111" when X = 146 AND Y = 15 else
"111111111111" when X = 147 AND Y = 15 else
"111111111111" when X = 148 AND Y = 15 else
"111111111111" when X = 149 AND Y = 15 else
"111111111111" when X = 150 AND Y = 15 else
"111111111111" when X = 151 AND Y = 15 else
"111111111111" when X = 152 AND Y = 15 else
"111111111111" when X = 153 AND Y = 15 else
"111111111111" when X = 154 AND Y = 15 else
"000000000000" when X = 155 AND Y = 15 else
"000000000000" when X = 156 AND Y = 15 else
"000000000000" when X = 157 AND Y = 15 else
"000000000000" when X = 158 AND Y = 15 else
"000000000000" when X = 159 AND Y = 15 else
"000000000000" when X = 160 AND Y = 15 else
"000000000000" when X = 161 AND Y = 15 else
"000000000000" when X = 162 AND Y = 15 else
"000000000000" when X = 163 AND Y = 15 else
"000000000000" when X = 164 AND Y = 15 else
"000000000000" when X = 165 AND Y = 15 else
"000000000000" when X = 166 AND Y = 15 else
"000000000000" when X = 167 AND Y = 15 else
"000000000000" when X = 168 AND Y = 15 else
"000000000000" when X = 169 AND Y = 15 else
"000000000000" when X = 170 AND Y = 15 else
"000000000000" when X = 171 AND Y = 15 else
"000000000000" when X = 172 AND Y = 15 else
"000000000000" when X = 173 AND Y = 15 else
"000000000000" when X = 174 AND Y = 15 else
"000000000000" when X = 175 AND Y = 15 else
"000000000000" when X = 176 AND Y = 15 else
"000000000000" when X = 177 AND Y = 15 else
"000000000000" when X = 178 AND Y = 15 else
"000000000000" when X = 179 AND Y = 15 else
"000000000000" when X = 180 AND Y = 15 else
"000000000000" when X = 181 AND Y = 15 else
"000000000000" when X = 182 AND Y = 15 else
"000000000000" when X = 183 AND Y = 15 else
"000000000000" when X = 184 AND Y = 15 else
"000000000000" when X = 185 AND Y = 15 else
"000000000000" when X = 186 AND Y = 15 else
"000000000000" when X = 187 AND Y = 15 else
"000000000000" when X = 188 AND Y = 15 else
"000000000000" when X = 189 AND Y = 15 else
"000000000000" when X = 190 AND Y = 15 else
"000000000000" when X = 191 AND Y = 15 else
"000000000000" when X = 192 AND Y = 15 else
"000000000000" when X = 193 AND Y = 15 else
"000000000000" when X = 194 AND Y = 15 else
"000000000000" when X = 195 AND Y = 15 else
"000000000000" when X = 196 AND Y = 15 else
"000000000000" when X = 197 AND Y = 15 else
"000000000000" when X = 198 AND Y = 15 else
"000000000000" when X = 199 AND Y = 15 else
"000000000000" when X = 200 AND Y = 15 else
"000000000000" when X = 201 AND Y = 15 else
"000000000000" when X = 202 AND Y = 15 else
"000000000000" when X = 203 AND Y = 15 else
"000000000000" when X = 204 AND Y = 15 else
"000000000000" when X = 205 AND Y = 15 else
"000000000000" when X = 206 AND Y = 15 else
"000000000000" when X = 207 AND Y = 15 else
"000000000000" when X = 208 AND Y = 15 else
"000000000000" when X = 209 AND Y = 15 else
"000000000000" when X = 210 AND Y = 15 else
"000000000000" when X = 211 AND Y = 15 else
"000000000000" when X = 212 AND Y = 15 else
"000000000000" when X = 213 AND Y = 15 else
"000000000000" when X = 214 AND Y = 15 else
"000000000000" when X = 215 AND Y = 15 else
"000000000000" when X = 216 AND Y = 15 else
"000000000000" when X = 217 AND Y = 15 else
"000000000000" when X = 218 AND Y = 15 else
"000000000000" when X = 219 AND Y = 15 else
"000000000000" when X = 220 AND Y = 15 else
"000000000000" when X = 221 AND Y = 15 else
"000000000000" when X = 222 AND Y = 15 else
"000000000000" when X = 223 AND Y = 15 else
"000000000000" when X = 224 AND Y = 15 else
"000000000000" when X = 225 AND Y = 15 else
"000000000000" when X = 226 AND Y = 15 else
"000000000000" when X = 227 AND Y = 15 else
"000000000000" when X = 228 AND Y = 15 else
"000000000000" when X = 229 AND Y = 15 else
"000000000000" when X = 230 AND Y = 15 else
"000000000000" when X = 231 AND Y = 15 else
"000000000000" when X = 232 AND Y = 15 else
"000000000000" when X = 233 AND Y = 15 else
"000000000000" when X = 234 AND Y = 15 else
"000000000000" when X = 235 AND Y = 15 else
"000000000000" when X = 236 AND Y = 15 else
"000000000000" when X = 237 AND Y = 15 else
"000000000000" when X = 238 AND Y = 15 else
"000000000000" when X = 239 AND Y = 15 else
"000000000000" when X = 240 AND Y = 15 else
"000000000000" when X = 241 AND Y = 15 else
"000000000000" when X = 242 AND Y = 15 else
"000000000000" when X = 243 AND Y = 15 else
"000000000000" when X = 244 AND Y = 15 else
"000000000000" when X = 245 AND Y = 15 else
"000000000000" when X = 246 AND Y = 15 else
"000000000000" when X = 247 AND Y = 15 else
"000000000000" when X = 248 AND Y = 15 else
"000000000000" when X = 249 AND Y = 15 else
"000000000000" when X = 250 AND Y = 15 else
"000000000000" when X = 251 AND Y = 15 else
"000000000000" when X = 252 AND Y = 15 else
"000000000000" when X = 253 AND Y = 15 else
"000000000000" when X = 254 AND Y = 15 else
"000000000000" when X = 255 AND Y = 15 else
"000000000000" when X = 256 AND Y = 15 else
"000000000000" when X = 257 AND Y = 15 else
"000000000000" when X = 258 AND Y = 15 else
"000000000000" when X = 259 AND Y = 15 else
"000000000000" when X = 260 AND Y = 15 else
"000000000000" when X = 261 AND Y = 15 else
"000000000000" when X = 262 AND Y = 15 else
"000000000000" when X = 263 AND Y = 15 else
"000000000000" when X = 264 AND Y = 15 else
"000000000000" when X = 265 AND Y = 15 else
"000000000000" when X = 266 AND Y = 15 else
"000000000000" when X = 267 AND Y = 15 else
"000000000000" when X = 268 AND Y = 15 else
"000000000000" when X = 269 AND Y = 15 else
"000000000000" when X = 270 AND Y = 15 else
"000000000000" when X = 271 AND Y = 15 else
"000000000000" when X = 272 AND Y = 15 else
"000000000000" when X = 273 AND Y = 15 else
"000000000000" when X = 274 AND Y = 15 else
"000000000000" when X = 275 AND Y = 15 else
"000000000000" when X = 276 AND Y = 15 else
"000000000000" when X = 277 AND Y = 15 else
"000000000000" when X = 278 AND Y = 15 else
"000000000000" when X = 279 AND Y = 15 else
"000000000000" when X = 280 AND Y = 15 else
"000000000000" when X = 281 AND Y = 15 else
"000000000000" when X = 282 AND Y = 15 else
"000000000000" when X = 283 AND Y = 15 else
"000000000000" when X = 284 AND Y = 15 else
"000000000000" when X = 285 AND Y = 15 else
"000000000000" when X = 286 AND Y = 15 else
"000000000000" when X = 287 AND Y = 15 else
"000000000000" when X = 288 AND Y = 15 else
"000000000000" when X = 289 AND Y = 15 else
"000000000000" when X = 290 AND Y = 15 else
"000000000000" when X = 291 AND Y = 15 else
"000000000000" when X = 292 AND Y = 15 else
"000000000000" when X = 293 AND Y = 15 else
"000000000000" when X = 294 AND Y = 15 else
"000000000000" when X = 295 AND Y = 15 else
"000000000000" when X = 296 AND Y = 15 else
"000000000000" when X = 297 AND Y = 15 else
"000000000000" when X = 298 AND Y = 15 else
"000000000000" when X = 299 AND Y = 15 else
"000000000000" when X = 300 AND Y = 15 else
"000000000000" when X = 301 AND Y = 15 else
"000000000000" when X = 302 AND Y = 15 else
"000000000000" when X = 303 AND Y = 15 else
"000000000000" when X = 304 AND Y = 15 else
"000000000000" when X = 305 AND Y = 15 else
"000000000000" when X = 306 AND Y = 15 else
"000000000000" when X = 307 AND Y = 15 else
"000000000000" when X = 308 AND Y = 15 else
"000000000000" when X = 309 AND Y = 15 else
"000000000000" when X = 310 AND Y = 15 else
"000000000000" when X = 311 AND Y = 15 else
"000000000000" when X = 312 AND Y = 15 else
"000000000000" when X = 313 AND Y = 15 else
"000000000000" when X = 314 AND Y = 15 else
"000000000000" when X = 315 AND Y = 15 else
"000000000000" when X = 316 AND Y = 15 else
"000000000000" when X = 317 AND Y = 15 else
"000000000000" when X = 318 AND Y = 15 else
"000000000000" when X = 319 AND Y = 15 else
"000000000000" when X = 320 AND Y = 15 else
"000000000000" when X = 321 AND Y = 15 else
"000000000000" when X = 322 AND Y = 15 else
"000000000000" when X = 323 AND Y = 15 else
"000000000000" when X = 324 AND Y = 15 else
"000000000000" when X = 0 AND Y = 16 else
"000000000000" when X = 1 AND Y = 16 else
"000000000000" when X = 2 AND Y = 16 else
"000000000000" when X = 3 AND Y = 16 else
"000000000000" when X = 4 AND Y = 16 else
"000000000000" when X = 5 AND Y = 16 else
"000000000000" when X = 6 AND Y = 16 else
"000000000000" when X = 7 AND Y = 16 else
"000000000000" when X = 8 AND Y = 16 else
"000000000000" when X = 9 AND Y = 16 else
"000000000000" when X = 10 AND Y = 16 else
"000000000000" when X = 11 AND Y = 16 else
"000000000000" when X = 12 AND Y = 16 else
"000000000000" when X = 13 AND Y = 16 else
"000000000000" when X = 14 AND Y = 16 else
"000000000000" when X = 15 AND Y = 16 else
"000000000000" when X = 16 AND Y = 16 else
"000000000000" when X = 17 AND Y = 16 else
"000000000000" when X = 18 AND Y = 16 else
"000000000000" when X = 19 AND Y = 16 else
"000000000000" when X = 20 AND Y = 16 else
"000000000000" when X = 21 AND Y = 16 else
"000000000000" when X = 22 AND Y = 16 else
"000000000000" when X = 23 AND Y = 16 else
"000000000000" when X = 24 AND Y = 16 else
"000000000000" when X = 25 AND Y = 16 else
"000000000000" when X = 26 AND Y = 16 else
"000000000000" when X = 27 AND Y = 16 else
"000000000000" when X = 28 AND Y = 16 else
"000000000000" when X = 29 AND Y = 16 else
"000000000000" when X = 30 AND Y = 16 else
"000000000000" when X = 31 AND Y = 16 else
"000000000000" when X = 32 AND Y = 16 else
"000000000000" when X = 33 AND Y = 16 else
"000000000000" when X = 34 AND Y = 16 else
"000000000000" when X = 35 AND Y = 16 else
"000000000000" when X = 36 AND Y = 16 else
"000000000000" when X = 37 AND Y = 16 else
"000000000000" when X = 38 AND Y = 16 else
"000000000000" when X = 39 AND Y = 16 else
"100010011101" when X = 40 AND Y = 16 else
"100010011101" when X = 41 AND Y = 16 else
"100010011101" when X = 42 AND Y = 16 else
"100010011101" when X = 43 AND Y = 16 else
"100010011101" when X = 44 AND Y = 16 else
"100010011101" when X = 45 AND Y = 16 else
"100010011101" when X = 46 AND Y = 16 else
"100010011101" when X = 47 AND Y = 16 else
"100010011101" when X = 48 AND Y = 16 else
"100010011101" when X = 49 AND Y = 16 else
"110111011111" when X = 50 AND Y = 16 else
"110111011111" when X = 51 AND Y = 16 else
"110111011111" when X = 52 AND Y = 16 else
"110111011111" when X = 53 AND Y = 16 else
"110111011111" when X = 54 AND Y = 16 else
"110111011111" when X = 55 AND Y = 16 else
"110111011111" when X = 56 AND Y = 16 else
"110111011111" when X = 57 AND Y = 16 else
"110111011111" when X = 58 AND Y = 16 else
"110111011111" when X = 59 AND Y = 16 else
"110111011111" when X = 60 AND Y = 16 else
"110111011111" when X = 61 AND Y = 16 else
"110111011111" when X = 62 AND Y = 16 else
"110111011111" when X = 63 AND Y = 16 else
"110111011111" when X = 64 AND Y = 16 else
"111111111111" when X = 65 AND Y = 16 else
"111111111111" when X = 66 AND Y = 16 else
"111111111111" when X = 67 AND Y = 16 else
"111111111111" when X = 68 AND Y = 16 else
"111111111111" when X = 69 AND Y = 16 else
"111111111111" when X = 70 AND Y = 16 else
"111111111111" when X = 71 AND Y = 16 else
"111111111111" when X = 72 AND Y = 16 else
"111111111111" when X = 73 AND Y = 16 else
"111111111111" when X = 74 AND Y = 16 else
"111111111111" when X = 75 AND Y = 16 else
"111111111111" when X = 76 AND Y = 16 else
"111111111111" when X = 77 AND Y = 16 else
"111111111111" when X = 78 AND Y = 16 else
"111111111111" when X = 79 AND Y = 16 else
"111111111111" when X = 80 AND Y = 16 else
"111111111111" when X = 81 AND Y = 16 else
"111111111111" when X = 82 AND Y = 16 else
"111111111111" when X = 83 AND Y = 16 else
"111111111111" when X = 84 AND Y = 16 else
"111111111111" when X = 85 AND Y = 16 else
"111111111111" when X = 86 AND Y = 16 else
"111111111111" when X = 87 AND Y = 16 else
"111111111111" when X = 88 AND Y = 16 else
"111111111111" when X = 89 AND Y = 16 else
"111111111111" when X = 90 AND Y = 16 else
"111111111111" when X = 91 AND Y = 16 else
"111111111111" when X = 92 AND Y = 16 else
"111111111111" when X = 93 AND Y = 16 else
"111111111111" when X = 94 AND Y = 16 else
"111111111111" when X = 95 AND Y = 16 else
"111111111111" when X = 96 AND Y = 16 else
"111111111111" when X = 97 AND Y = 16 else
"111111111111" when X = 98 AND Y = 16 else
"111111111111" when X = 99 AND Y = 16 else
"111111111111" when X = 100 AND Y = 16 else
"111111111111" when X = 101 AND Y = 16 else
"111111111111" when X = 102 AND Y = 16 else
"111111111111" when X = 103 AND Y = 16 else
"111111111111" when X = 104 AND Y = 16 else
"111111111111" when X = 105 AND Y = 16 else
"111111111111" when X = 106 AND Y = 16 else
"111111111111" when X = 107 AND Y = 16 else
"111111111111" when X = 108 AND Y = 16 else
"111111111111" when X = 109 AND Y = 16 else
"111111111111" when X = 110 AND Y = 16 else
"111111111111" when X = 111 AND Y = 16 else
"111111111111" when X = 112 AND Y = 16 else
"111111111111" when X = 113 AND Y = 16 else
"111111111111" when X = 114 AND Y = 16 else
"111111111111" when X = 115 AND Y = 16 else
"111111111111" when X = 116 AND Y = 16 else
"111111111111" when X = 117 AND Y = 16 else
"111111111111" when X = 118 AND Y = 16 else
"111111111111" when X = 119 AND Y = 16 else
"111111111111" when X = 120 AND Y = 16 else
"111111111111" when X = 121 AND Y = 16 else
"111111111111" when X = 122 AND Y = 16 else
"111111111111" when X = 123 AND Y = 16 else
"111111111111" when X = 124 AND Y = 16 else
"111111111111" when X = 125 AND Y = 16 else
"111111111111" when X = 126 AND Y = 16 else
"111111111111" when X = 127 AND Y = 16 else
"111111111111" when X = 128 AND Y = 16 else
"111111111111" when X = 129 AND Y = 16 else
"111111111111" when X = 130 AND Y = 16 else
"111111111111" when X = 131 AND Y = 16 else
"111111111111" when X = 132 AND Y = 16 else
"111111111111" when X = 133 AND Y = 16 else
"111111111111" when X = 134 AND Y = 16 else
"111111111111" when X = 135 AND Y = 16 else
"111111111111" when X = 136 AND Y = 16 else
"111111111111" when X = 137 AND Y = 16 else
"111111111111" when X = 138 AND Y = 16 else
"111111111111" when X = 139 AND Y = 16 else
"111111111111" when X = 140 AND Y = 16 else
"111111111111" when X = 141 AND Y = 16 else
"111111111111" when X = 142 AND Y = 16 else
"111111111111" when X = 143 AND Y = 16 else
"111111111111" when X = 144 AND Y = 16 else
"111111111111" when X = 145 AND Y = 16 else
"111111111111" when X = 146 AND Y = 16 else
"111111111111" when X = 147 AND Y = 16 else
"111111111111" when X = 148 AND Y = 16 else
"111111111111" when X = 149 AND Y = 16 else
"111111111111" when X = 150 AND Y = 16 else
"111111111111" when X = 151 AND Y = 16 else
"111111111111" when X = 152 AND Y = 16 else
"111111111111" when X = 153 AND Y = 16 else
"111111111111" when X = 154 AND Y = 16 else
"000000000000" when X = 155 AND Y = 16 else
"000000000000" when X = 156 AND Y = 16 else
"000000000000" when X = 157 AND Y = 16 else
"000000000000" when X = 158 AND Y = 16 else
"000000000000" when X = 159 AND Y = 16 else
"000000000000" when X = 160 AND Y = 16 else
"000000000000" when X = 161 AND Y = 16 else
"000000000000" when X = 162 AND Y = 16 else
"000000000000" when X = 163 AND Y = 16 else
"000000000000" when X = 164 AND Y = 16 else
"000000000000" when X = 165 AND Y = 16 else
"000000000000" when X = 166 AND Y = 16 else
"000000000000" when X = 167 AND Y = 16 else
"000000000000" when X = 168 AND Y = 16 else
"000000000000" when X = 169 AND Y = 16 else
"000000000000" when X = 170 AND Y = 16 else
"000000000000" when X = 171 AND Y = 16 else
"000000000000" when X = 172 AND Y = 16 else
"000000000000" when X = 173 AND Y = 16 else
"000000000000" when X = 174 AND Y = 16 else
"000000000000" when X = 175 AND Y = 16 else
"000000000000" when X = 176 AND Y = 16 else
"000000000000" when X = 177 AND Y = 16 else
"000000000000" when X = 178 AND Y = 16 else
"000000000000" when X = 179 AND Y = 16 else
"000000000000" when X = 180 AND Y = 16 else
"000000000000" when X = 181 AND Y = 16 else
"000000000000" when X = 182 AND Y = 16 else
"000000000000" when X = 183 AND Y = 16 else
"000000000000" when X = 184 AND Y = 16 else
"000000000000" when X = 185 AND Y = 16 else
"000000000000" when X = 186 AND Y = 16 else
"000000000000" when X = 187 AND Y = 16 else
"000000000000" when X = 188 AND Y = 16 else
"000000000000" when X = 189 AND Y = 16 else
"000000000000" when X = 190 AND Y = 16 else
"000000000000" when X = 191 AND Y = 16 else
"000000000000" when X = 192 AND Y = 16 else
"000000000000" when X = 193 AND Y = 16 else
"000000000000" when X = 194 AND Y = 16 else
"000000000000" when X = 195 AND Y = 16 else
"000000000000" when X = 196 AND Y = 16 else
"000000000000" when X = 197 AND Y = 16 else
"000000000000" when X = 198 AND Y = 16 else
"000000000000" when X = 199 AND Y = 16 else
"000000000000" when X = 200 AND Y = 16 else
"000000000000" when X = 201 AND Y = 16 else
"000000000000" when X = 202 AND Y = 16 else
"000000000000" when X = 203 AND Y = 16 else
"000000000000" when X = 204 AND Y = 16 else
"000000000000" when X = 205 AND Y = 16 else
"000000000000" when X = 206 AND Y = 16 else
"000000000000" when X = 207 AND Y = 16 else
"000000000000" when X = 208 AND Y = 16 else
"000000000000" when X = 209 AND Y = 16 else
"000000000000" when X = 210 AND Y = 16 else
"000000000000" when X = 211 AND Y = 16 else
"000000000000" when X = 212 AND Y = 16 else
"000000000000" when X = 213 AND Y = 16 else
"000000000000" when X = 214 AND Y = 16 else
"000000000000" when X = 215 AND Y = 16 else
"000000000000" when X = 216 AND Y = 16 else
"000000000000" when X = 217 AND Y = 16 else
"000000000000" when X = 218 AND Y = 16 else
"000000000000" when X = 219 AND Y = 16 else
"000000000000" when X = 220 AND Y = 16 else
"000000000000" when X = 221 AND Y = 16 else
"000000000000" when X = 222 AND Y = 16 else
"000000000000" when X = 223 AND Y = 16 else
"000000000000" when X = 224 AND Y = 16 else
"000000000000" when X = 225 AND Y = 16 else
"000000000000" when X = 226 AND Y = 16 else
"000000000000" when X = 227 AND Y = 16 else
"000000000000" when X = 228 AND Y = 16 else
"000000000000" when X = 229 AND Y = 16 else
"000000000000" when X = 230 AND Y = 16 else
"000000000000" when X = 231 AND Y = 16 else
"000000000000" when X = 232 AND Y = 16 else
"000000000000" when X = 233 AND Y = 16 else
"000000000000" when X = 234 AND Y = 16 else
"000000000000" when X = 235 AND Y = 16 else
"000000000000" when X = 236 AND Y = 16 else
"000000000000" when X = 237 AND Y = 16 else
"000000000000" when X = 238 AND Y = 16 else
"000000000000" when X = 239 AND Y = 16 else
"000000000000" when X = 240 AND Y = 16 else
"000000000000" when X = 241 AND Y = 16 else
"000000000000" when X = 242 AND Y = 16 else
"000000000000" when X = 243 AND Y = 16 else
"000000000000" when X = 244 AND Y = 16 else
"000000000000" when X = 245 AND Y = 16 else
"000000000000" when X = 246 AND Y = 16 else
"000000000000" when X = 247 AND Y = 16 else
"000000000000" when X = 248 AND Y = 16 else
"000000000000" when X = 249 AND Y = 16 else
"000000000000" when X = 250 AND Y = 16 else
"000000000000" when X = 251 AND Y = 16 else
"000000000000" when X = 252 AND Y = 16 else
"000000000000" when X = 253 AND Y = 16 else
"000000000000" when X = 254 AND Y = 16 else
"000000000000" when X = 255 AND Y = 16 else
"000000000000" when X = 256 AND Y = 16 else
"000000000000" when X = 257 AND Y = 16 else
"000000000000" when X = 258 AND Y = 16 else
"000000000000" when X = 259 AND Y = 16 else
"000000000000" when X = 260 AND Y = 16 else
"000000000000" when X = 261 AND Y = 16 else
"000000000000" when X = 262 AND Y = 16 else
"000000000000" when X = 263 AND Y = 16 else
"000000000000" when X = 264 AND Y = 16 else
"000000000000" when X = 265 AND Y = 16 else
"000000000000" when X = 266 AND Y = 16 else
"000000000000" when X = 267 AND Y = 16 else
"000000000000" when X = 268 AND Y = 16 else
"000000000000" when X = 269 AND Y = 16 else
"000000000000" when X = 270 AND Y = 16 else
"000000000000" when X = 271 AND Y = 16 else
"000000000000" when X = 272 AND Y = 16 else
"000000000000" when X = 273 AND Y = 16 else
"000000000000" when X = 274 AND Y = 16 else
"000000000000" when X = 275 AND Y = 16 else
"000000000000" when X = 276 AND Y = 16 else
"000000000000" when X = 277 AND Y = 16 else
"000000000000" when X = 278 AND Y = 16 else
"000000000000" when X = 279 AND Y = 16 else
"000000000000" when X = 280 AND Y = 16 else
"000000000000" when X = 281 AND Y = 16 else
"000000000000" when X = 282 AND Y = 16 else
"000000000000" when X = 283 AND Y = 16 else
"000000000000" when X = 284 AND Y = 16 else
"000000000000" when X = 285 AND Y = 16 else
"000000000000" when X = 286 AND Y = 16 else
"000000000000" when X = 287 AND Y = 16 else
"000000000000" when X = 288 AND Y = 16 else
"000000000000" when X = 289 AND Y = 16 else
"000000000000" when X = 290 AND Y = 16 else
"000000000000" when X = 291 AND Y = 16 else
"000000000000" when X = 292 AND Y = 16 else
"000000000000" when X = 293 AND Y = 16 else
"000000000000" when X = 294 AND Y = 16 else
"000000000000" when X = 295 AND Y = 16 else
"000000000000" when X = 296 AND Y = 16 else
"000000000000" when X = 297 AND Y = 16 else
"000000000000" when X = 298 AND Y = 16 else
"000000000000" when X = 299 AND Y = 16 else
"000000000000" when X = 300 AND Y = 16 else
"000000000000" when X = 301 AND Y = 16 else
"000000000000" when X = 302 AND Y = 16 else
"000000000000" when X = 303 AND Y = 16 else
"000000000000" when X = 304 AND Y = 16 else
"000000000000" when X = 305 AND Y = 16 else
"000000000000" when X = 306 AND Y = 16 else
"000000000000" when X = 307 AND Y = 16 else
"000000000000" when X = 308 AND Y = 16 else
"000000000000" when X = 309 AND Y = 16 else
"000000000000" when X = 310 AND Y = 16 else
"000000000000" when X = 311 AND Y = 16 else
"000000000000" when X = 312 AND Y = 16 else
"000000000000" when X = 313 AND Y = 16 else
"000000000000" when X = 314 AND Y = 16 else
"000000000000" when X = 315 AND Y = 16 else
"000000000000" when X = 316 AND Y = 16 else
"000000000000" when X = 317 AND Y = 16 else
"000000000000" when X = 318 AND Y = 16 else
"000000000000" when X = 319 AND Y = 16 else
"000000000000" when X = 320 AND Y = 16 else
"000000000000" when X = 321 AND Y = 16 else
"000000000000" when X = 322 AND Y = 16 else
"000000000000" when X = 323 AND Y = 16 else
"000000000000" when X = 324 AND Y = 16 else
"000000000000" when X = 0 AND Y = 17 else
"000000000000" when X = 1 AND Y = 17 else
"000000000000" when X = 2 AND Y = 17 else
"000000000000" when X = 3 AND Y = 17 else
"000000000000" when X = 4 AND Y = 17 else
"000000000000" when X = 5 AND Y = 17 else
"000000000000" when X = 6 AND Y = 17 else
"000000000000" when X = 7 AND Y = 17 else
"000000000000" when X = 8 AND Y = 17 else
"000000000000" when X = 9 AND Y = 17 else
"000000000000" when X = 10 AND Y = 17 else
"000000000000" when X = 11 AND Y = 17 else
"000000000000" when X = 12 AND Y = 17 else
"000000000000" when X = 13 AND Y = 17 else
"000000000000" when X = 14 AND Y = 17 else
"000000000000" when X = 15 AND Y = 17 else
"000000000000" when X = 16 AND Y = 17 else
"000000000000" when X = 17 AND Y = 17 else
"000000000000" when X = 18 AND Y = 17 else
"000000000000" when X = 19 AND Y = 17 else
"000000000000" when X = 20 AND Y = 17 else
"000000000000" when X = 21 AND Y = 17 else
"000000000000" when X = 22 AND Y = 17 else
"000000000000" when X = 23 AND Y = 17 else
"000000000000" when X = 24 AND Y = 17 else
"000000000000" when X = 25 AND Y = 17 else
"000000000000" when X = 26 AND Y = 17 else
"000000000000" when X = 27 AND Y = 17 else
"000000000000" when X = 28 AND Y = 17 else
"000000000000" when X = 29 AND Y = 17 else
"000000000000" when X = 30 AND Y = 17 else
"000000000000" when X = 31 AND Y = 17 else
"000000000000" when X = 32 AND Y = 17 else
"000000000000" when X = 33 AND Y = 17 else
"000000000000" when X = 34 AND Y = 17 else
"000000000000" when X = 35 AND Y = 17 else
"000000000000" when X = 36 AND Y = 17 else
"000000000000" when X = 37 AND Y = 17 else
"000000000000" when X = 38 AND Y = 17 else
"000000000000" when X = 39 AND Y = 17 else
"100010011101" when X = 40 AND Y = 17 else
"100010011101" when X = 41 AND Y = 17 else
"100010011101" when X = 42 AND Y = 17 else
"100010011101" when X = 43 AND Y = 17 else
"100010011101" when X = 44 AND Y = 17 else
"100010011101" when X = 45 AND Y = 17 else
"100010011101" when X = 46 AND Y = 17 else
"100010011101" when X = 47 AND Y = 17 else
"100010011101" when X = 48 AND Y = 17 else
"100010011101" when X = 49 AND Y = 17 else
"110111011111" when X = 50 AND Y = 17 else
"110111011111" when X = 51 AND Y = 17 else
"110111011111" when X = 52 AND Y = 17 else
"110111011111" when X = 53 AND Y = 17 else
"110111011111" when X = 54 AND Y = 17 else
"110111011111" when X = 55 AND Y = 17 else
"110111011111" when X = 56 AND Y = 17 else
"110111011111" when X = 57 AND Y = 17 else
"110111011111" when X = 58 AND Y = 17 else
"110111011111" when X = 59 AND Y = 17 else
"110111011111" when X = 60 AND Y = 17 else
"110111011111" when X = 61 AND Y = 17 else
"110111011111" when X = 62 AND Y = 17 else
"110111011111" when X = 63 AND Y = 17 else
"110111011111" when X = 64 AND Y = 17 else
"111111111111" when X = 65 AND Y = 17 else
"111111111111" when X = 66 AND Y = 17 else
"111111111111" when X = 67 AND Y = 17 else
"111111111111" when X = 68 AND Y = 17 else
"111111111111" when X = 69 AND Y = 17 else
"111111111111" when X = 70 AND Y = 17 else
"111111111111" when X = 71 AND Y = 17 else
"111111111111" when X = 72 AND Y = 17 else
"111111111111" when X = 73 AND Y = 17 else
"111111111111" when X = 74 AND Y = 17 else
"111111111111" when X = 75 AND Y = 17 else
"111111111111" when X = 76 AND Y = 17 else
"111111111111" when X = 77 AND Y = 17 else
"111111111111" when X = 78 AND Y = 17 else
"111111111111" when X = 79 AND Y = 17 else
"111111111111" when X = 80 AND Y = 17 else
"111111111111" when X = 81 AND Y = 17 else
"111111111111" when X = 82 AND Y = 17 else
"111111111111" when X = 83 AND Y = 17 else
"111111111111" when X = 84 AND Y = 17 else
"111111111111" when X = 85 AND Y = 17 else
"111111111111" when X = 86 AND Y = 17 else
"111111111111" when X = 87 AND Y = 17 else
"111111111111" when X = 88 AND Y = 17 else
"111111111111" when X = 89 AND Y = 17 else
"111111111111" when X = 90 AND Y = 17 else
"111111111111" when X = 91 AND Y = 17 else
"111111111111" when X = 92 AND Y = 17 else
"111111111111" when X = 93 AND Y = 17 else
"111111111111" when X = 94 AND Y = 17 else
"111111111111" when X = 95 AND Y = 17 else
"111111111111" when X = 96 AND Y = 17 else
"111111111111" when X = 97 AND Y = 17 else
"111111111111" when X = 98 AND Y = 17 else
"111111111111" when X = 99 AND Y = 17 else
"111111111111" when X = 100 AND Y = 17 else
"111111111111" when X = 101 AND Y = 17 else
"111111111111" when X = 102 AND Y = 17 else
"111111111111" when X = 103 AND Y = 17 else
"111111111111" when X = 104 AND Y = 17 else
"111111111111" when X = 105 AND Y = 17 else
"111111111111" when X = 106 AND Y = 17 else
"111111111111" when X = 107 AND Y = 17 else
"111111111111" when X = 108 AND Y = 17 else
"111111111111" when X = 109 AND Y = 17 else
"111111111111" when X = 110 AND Y = 17 else
"111111111111" when X = 111 AND Y = 17 else
"111111111111" when X = 112 AND Y = 17 else
"111111111111" when X = 113 AND Y = 17 else
"111111111111" when X = 114 AND Y = 17 else
"111111111111" when X = 115 AND Y = 17 else
"111111111111" when X = 116 AND Y = 17 else
"111111111111" when X = 117 AND Y = 17 else
"111111111111" when X = 118 AND Y = 17 else
"111111111111" when X = 119 AND Y = 17 else
"111111111111" when X = 120 AND Y = 17 else
"111111111111" when X = 121 AND Y = 17 else
"111111111111" when X = 122 AND Y = 17 else
"111111111111" when X = 123 AND Y = 17 else
"111111111111" when X = 124 AND Y = 17 else
"111111111111" when X = 125 AND Y = 17 else
"111111111111" when X = 126 AND Y = 17 else
"111111111111" when X = 127 AND Y = 17 else
"111111111111" when X = 128 AND Y = 17 else
"111111111111" when X = 129 AND Y = 17 else
"111111111111" when X = 130 AND Y = 17 else
"111111111111" when X = 131 AND Y = 17 else
"111111111111" when X = 132 AND Y = 17 else
"111111111111" when X = 133 AND Y = 17 else
"111111111111" when X = 134 AND Y = 17 else
"111111111111" when X = 135 AND Y = 17 else
"111111111111" when X = 136 AND Y = 17 else
"111111111111" when X = 137 AND Y = 17 else
"111111111111" when X = 138 AND Y = 17 else
"111111111111" when X = 139 AND Y = 17 else
"111111111111" when X = 140 AND Y = 17 else
"111111111111" when X = 141 AND Y = 17 else
"111111111111" when X = 142 AND Y = 17 else
"111111111111" when X = 143 AND Y = 17 else
"111111111111" when X = 144 AND Y = 17 else
"111111111111" when X = 145 AND Y = 17 else
"111111111111" when X = 146 AND Y = 17 else
"111111111111" when X = 147 AND Y = 17 else
"111111111111" when X = 148 AND Y = 17 else
"111111111111" when X = 149 AND Y = 17 else
"111111111111" when X = 150 AND Y = 17 else
"111111111111" when X = 151 AND Y = 17 else
"111111111111" when X = 152 AND Y = 17 else
"111111111111" when X = 153 AND Y = 17 else
"111111111111" when X = 154 AND Y = 17 else
"000000000000" when X = 155 AND Y = 17 else
"000000000000" when X = 156 AND Y = 17 else
"000000000000" when X = 157 AND Y = 17 else
"000000000000" when X = 158 AND Y = 17 else
"000000000000" when X = 159 AND Y = 17 else
"000000000000" when X = 160 AND Y = 17 else
"000000000000" when X = 161 AND Y = 17 else
"000000000000" when X = 162 AND Y = 17 else
"000000000000" when X = 163 AND Y = 17 else
"000000000000" when X = 164 AND Y = 17 else
"000000000000" when X = 165 AND Y = 17 else
"000000000000" when X = 166 AND Y = 17 else
"000000000000" when X = 167 AND Y = 17 else
"000000000000" when X = 168 AND Y = 17 else
"000000000000" when X = 169 AND Y = 17 else
"000000000000" when X = 170 AND Y = 17 else
"000000000000" when X = 171 AND Y = 17 else
"000000000000" when X = 172 AND Y = 17 else
"000000000000" when X = 173 AND Y = 17 else
"000000000000" when X = 174 AND Y = 17 else
"000000000000" when X = 175 AND Y = 17 else
"000000000000" when X = 176 AND Y = 17 else
"000000000000" when X = 177 AND Y = 17 else
"000000000000" when X = 178 AND Y = 17 else
"000000000000" when X = 179 AND Y = 17 else
"000000000000" when X = 180 AND Y = 17 else
"000000000000" when X = 181 AND Y = 17 else
"000000000000" when X = 182 AND Y = 17 else
"000000000000" when X = 183 AND Y = 17 else
"000000000000" when X = 184 AND Y = 17 else
"000000000000" when X = 185 AND Y = 17 else
"000000000000" when X = 186 AND Y = 17 else
"000000000000" when X = 187 AND Y = 17 else
"000000000000" when X = 188 AND Y = 17 else
"000000000000" when X = 189 AND Y = 17 else
"000000000000" when X = 190 AND Y = 17 else
"000000000000" when X = 191 AND Y = 17 else
"000000000000" when X = 192 AND Y = 17 else
"000000000000" when X = 193 AND Y = 17 else
"000000000000" when X = 194 AND Y = 17 else
"000000000000" when X = 195 AND Y = 17 else
"000000000000" when X = 196 AND Y = 17 else
"000000000000" when X = 197 AND Y = 17 else
"000000000000" when X = 198 AND Y = 17 else
"000000000000" when X = 199 AND Y = 17 else
"000000000000" when X = 200 AND Y = 17 else
"000000000000" when X = 201 AND Y = 17 else
"000000000000" when X = 202 AND Y = 17 else
"000000000000" when X = 203 AND Y = 17 else
"000000000000" when X = 204 AND Y = 17 else
"000000000000" when X = 205 AND Y = 17 else
"000000000000" when X = 206 AND Y = 17 else
"000000000000" when X = 207 AND Y = 17 else
"000000000000" when X = 208 AND Y = 17 else
"000000000000" when X = 209 AND Y = 17 else
"000000000000" when X = 210 AND Y = 17 else
"000000000000" when X = 211 AND Y = 17 else
"000000000000" when X = 212 AND Y = 17 else
"000000000000" when X = 213 AND Y = 17 else
"000000000000" when X = 214 AND Y = 17 else
"000000000000" when X = 215 AND Y = 17 else
"000000000000" when X = 216 AND Y = 17 else
"000000000000" when X = 217 AND Y = 17 else
"000000000000" when X = 218 AND Y = 17 else
"000000000000" when X = 219 AND Y = 17 else
"000000000000" when X = 220 AND Y = 17 else
"000000000000" when X = 221 AND Y = 17 else
"000000000000" when X = 222 AND Y = 17 else
"000000000000" when X = 223 AND Y = 17 else
"000000000000" when X = 224 AND Y = 17 else
"000000000000" when X = 225 AND Y = 17 else
"000000000000" when X = 226 AND Y = 17 else
"000000000000" when X = 227 AND Y = 17 else
"000000000000" when X = 228 AND Y = 17 else
"000000000000" when X = 229 AND Y = 17 else
"000000000000" when X = 230 AND Y = 17 else
"000000000000" when X = 231 AND Y = 17 else
"000000000000" when X = 232 AND Y = 17 else
"000000000000" when X = 233 AND Y = 17 else
"000000000000" when X = 234 AND Y = 17 else
"000000000000" when X = 235 AND Y = 17 else
"000000000000" when X = 236 AND Y = 17 else
"000000000000" when X = 237 AND Y = 17 else
"000000000000" when X = 238 AND Y = 17 else
"000000000000" when X = 239 AND Y = 17 else
"000000000000" when X = 240 AND Y = 17 else
"000000000000" when X = 241 AND Y = 17 else
"000000000000" when X = 242 AND Y = 17 else
"000000000000" when X = 243 AND Y = 17 else
"000000000000" when X = 244 AND Y = 17 else
"000000000000" when X = 245 AND Y = 17 else
"000000000000" when X = 246 AND Y = 17 else
"000000000000" when X = 247 AND Y = 17 else
"000000000000" when X = 248 AND Y = 17 else
"000000000000" when X = 249 AND Y = 17 else
"000000000000" when X = 250 AND Y = 17 else
"000000000000" when X = 251 AND Y = 17 else
"000000000000" when X = 252 AND Y = 17 else
"000000000000" when X = 253 AND Y = 17 else
"000000000000" when X = 254 AND Y = 17 else
"000000000000" when X = 255 AND Y = 17 else
"000000000000" when X = 256 AND Y = 17 else
"000000000000" when X = 257 AND Y = 17 else
"000000000000" when X = 258 AND Y = 17 else
"000000000000" when X = 259 AND Y = 17 else
"000000000000" when X = 260 AND Y = 17 else
"000000000000" when X = 261 AND Y = 17 else
"000000000000" when X = 262 AND Y = 17 else
"000000000000" when X = 263 AND Y = 17 else
"000000000000" when X = 264 AND Y = 17 else
"000000000000" when X = 265 AND Y = 17 else
"000000000000" when X = 266 AND Y = 17 else
"000000000000" when X = 267 AND Y = 17 else
"000000000000" when X = 268 AND Y = 17 else
"000000000000" when X = 269 AND Y = 17 else
"000000000000" when X = 270 AND Y = 17 else
"000000000000" when X = 271 AND Y = 17 else
"000000000000" when X = 272 AND Y = 17 else
"000000000000" when X = 273 AND Y = 17 else
"000000000000" when X = 274 AND Y = 17 else
"000000000000" when X = 275 AND Y = 17 else
"000000000000" when X = 276 AND Y = 17 else
"000000000000" when X = 277 AND Y = 17 else
"000000000000" when X = 278 AND Y = 17 else
"000000000000" when X = 279 AND Y = 17 else
"000000000000" when X = 280 AND Y = 17 else
"000000000000" when X = 281 AND Y = 17 else
"000000000000" when X = 282 AND Y = 17 else
"000000000000" when X = 283 AND Y = 17 else
"000000000000" when X = 284 AND Y = 17 else
"000000000000" when X = 285 AND Y = 17 else
"000000000000" when X = 286 AND Y = 17 else
"000000000000" when X = 287 AND Y = 17 else
"000000000000" when X = 288 AND Y = 17 else
"000000000000" when X = 289 AND Y = 17 else
"000000000000" when X = 290 AND Y = 17 else
"000000000000" when X = 291 AND Y = 17 else
"000000000000" when X = 292 AND Y = 17 else
"000000000000" when X = 293 AND Y = 17 else
"000000000000" when X = 294 AND Y = 17 else
"000000000000" when X = 295 AND Y = 17 else
"000000000000" when X = 296 AND Y = 17 else
"000000000000" when X = 297 AND Y = 17 else
"000000000000" when X = 298 AND Y = 17 else
"000000000000" when X = 299 AND Y = 17 else
"000000000000" when X = 300 AND Y = 17 else
"000000000000" when X = 301 AND Y = 17 else
"000000000000" when X = 302 AND Y = 17 else
"000000000000" when X = 303 AND Y = 17 else
"000000000000" when X = 304 AND Y = 17 else
"000000000000" when X = 305 AND Y = 17 else
"000000000000" when X = 306 AND Y = 17 else
"000000000000" when X = 307 AND Y = 17 else
"000000000000" when X = 308 AND Y = 17 else
"000000000000" when X = 309 AND Y = 17 else
"000000000000" when X = 310 AND Y = 17 else
"000000000000" when X = 311 AND Y = 17 else
"000000000000" when X = 312 AND Y = 17 else
"000000000000" when X = 313 AND Y = 17 else
"000000000000" when X = 314 AND Y = 17 else
"000000000000" when X = 315 AND Y = 17 else
"000000000000" when X = 316 AND Y = 17 else
"000000000000" when X = 317 AND Y = 17 else
"000000000000" when X = 318 AND Y = 17 else
"000000000000" when X = 319 AND Y = 17 else
"000000000000" when X = 320 AND Y = 17 else
"000000000000" when X = 321 AND Y = 17 else
"000000000000" when X = 322 AND Y = 17 else
"000000000000" when X = 323 AND Y = 17 else
"000000000000" when X = 324 AND Y = 17 else
"000000000000" when X = 0 AND Y = 18 else
"000000000000" when X = 1 AND Y = 18 else
"000000000000" when X = 2 AND Y = 18 else
"000000000000" when X = 3 AND Y = 18 else
"000000000000" when X = 4 AND Y = 18 else
"000000000000" when X = 5 AND Y = 18 else
"000000000000" when X = 6 AND Y = 18 else
"000000000000" when X = 7 AND Y = 18 else
"000000000000" when X = 8 AND Y = 18 else
"000000000000" when X = 9 AND Y = 18 else
"000000000000" when X = 10 AND Y = 18 else
"000000000000" when X = 11 AND Y = 18 else
"000000000000" when X = 12 AND Y = 18 else
"000000000000" when X = 13 AND Y = 18 else
"000000000000" when X = 14 AND Y = 18 else
"000000000000" when X = 15 AND Y = 18 else
"000000000000" when X = 16 AND Y = 18 else
"000000000000" when X = 17 AND Y = 18 else
"000000000000" when X = 18 AND Y = 18 else
"000000000000" when X = 19 AND Y = 18 else
"000000000000" when X = 20 AND Y = 18 else
"000000000000" when X = 21 AND Y = 18 else
"000000000000" when X = 22 AND Y = 18 else
"000000000000" when X = 23 AND Y = 18 else
"000000000000" when X = 24 AND Y = 18 else
"000000000000" when X = 25 AND Y = 18 else
"000000000000" when X = 26 AND Y = 18 else
"000000000000" when X = 27 AND Y = 18 else
"000000000000" when X = 28 AND Y = 18 else
"000000000000" when X = 29 AND Y = 18 else
"000000000000" when X = 30 AND Y = 18 else
"000000000000" when X = 31 AND Y = 18 else
"000000000000" when X = 32 AND Y = 18 else
"000000000000" when X = 33 AND Y = 18 else
"000000000000" when X = 34 AND Y = 18 else
"000000000000" when X = 35 AND Y = 18 else
"000000000000" when X = 36 AND Y = 18 else
"000000000000" when X = 37 AND Y = 18 else
"000000000000" when X = 38 AND Y = 18 else
"000000000000" when X = 39 AND Y = 18 else
"100010011101" when X = 40 AND Y = 18 else
"100010011101" when X = 41 AND Y = 18 else
"100010011101" when X = 42 AND Y = 18 else
"100010011101" when X = 43 AND Y = 18 else
"100010011101" when X = 44 AND Y = 18 else
"100010011101" when X = 45 AND Y = 18 else
"100010011101" when X = 46 AND Y = 18 else
"100010011101" when X = 47 AND Y = 18 else
"100010011101" when X = 48 AND Y = 18 else
"100010011101" when X = 49 AND Y = 18 else
"110111011111" when X = 50 AND Y = 18 else
"110111011111" when X = 51 AND Y = 18 else
"110111011111" when X = 52 AND Y = 18 else
"110111011111" when X = 53 AND Y = 18 else
"110111011111" when X = 54 AND Y = 18 else
"110111011111" when X = 55 AND Y = 18 else
"110111011111" when X = 56 AND Y = 18 else
"110111011111" when X = 57 AND Y = 18 else
"110111011111" when X = 58 AND Y = 18 else
"110111011111" when X = 59 AND Y = 18 else
"110111011111" when X = 60 AND Y = 18 else
"110111011111" when X = 61 AND Y = 18 else
"110111011111" when X = 62 AND Y = 18 else
"110111011111" when X = 63 AND Y = 18 else
"110111011111" when X = 64 AND Y = 18 else
"111111111111" when X = 65 AND Y = 18 else
"111111111111" when X = 66 AND Y = 18 else
"111111111111" when X = 67 AND Y = 18 else
"111111111111" when X = 68 AND Y = 18 else
"111111111111" when X = 69 AND Y = 18 else
"111111111111" when X = 70 AND Y = 18 else
"111111111111" when X = 71 AND Y = 18 else
"111111111111" when X = 72 AND Y = 18 else
"111111111111" when X = 73 AND Y = 18 else
"111111111111" when X = 74 AND Y = 18 else
"111111111111" when X = 75 AND Y = 18 else
"111111111111" when X = 76 AND Y = 18 else
"111111111111" when X = 77 AND Y = 18 else
"111111111111" when X = 78 AND Y = 18 else
"111111111111" when X = 79 AND Y = 18 else
"111111111111" when X = 80 AND Y = 18 else
"111111111111" when X = 81 AND Y = 18 else
"111111111111" when X = 82 AND Y = 18 else
"111111111111" when X = 83 AND Y = 18 else
"111111111111" when X = 84 AND Y = 18 else
"111111111111" when X = 85 AND Y = 18 else
"111111111111" when X = 86 AND Y = 18 else
"111111111111" when X = 87 AND Y = 18 else
"111111111111" when X = 88 AND Y = 18 else
"111111111111" when X = 89 AND Y = 18 else
"111111111111" when X = 90 AND Y = 18 else
"111111111111" when X = 91 AND Y = 18 else
"111111111111" when X = 92 AND Y = 18 else
"111111111111" when X = 93 AND Y = 18 else
"111111111111" when X = 94 AND Y = 18 else
"111111111111" when X = 95 AND Y = 18 else
"111111111111" when X = 96 AND Y = 18 else
"111111111111" when X = 97 AND Y = 18 else
"111111111111" when X = 98 AND Y = 18 else
"111111111111" when X = 99 AND Y = 18 else
"111111111111" when X = 100 AND Y = 18 else
"111111111111" when X = 101 AND Y = 18 else
"111111111111" when X = 102 AND Y = 18 else
"111111111111" when X = 103 AND Y = 18 else
"111111111111" when X = 104 AND Y = 18 else
"111111111111" when X = 105 AND Y = 18 else
"111111111111" when X = 106 AND Y = 18 else
"111111111111" when X = 107 AND Y = 18 else
"111111111111" when X = 108 AND Y = 18 else
"111111111111" when X = 109 AND Y = 18 else
"111111111111" when X = 110 AND Y = 18 else
"111111111111" when X = 111 AND Y = 18 else
"111111111111" when X = 112 AND Y = 18 else
"111111111111" when X = 113 AND Y = 18 else
"111111111111" when X = 114 AND Y = 18 else
"111111111111" when X = 115 AND Y = 18 else
"111111111111" when X = 116 AND Y = 18 else
"111111111111" when X = 117 AND Y = 18 else
"111111111111" when X = 118 AND Y = 18 else
"111111111111" when X = 119 AND Y = 18 else
"111111111111" when X = 120 AND Y = 18 else
"111111111111" when X = 121 AND Y = 18 else
"111111111111" when X = 122 AND Y = 18 else
"111111111111" when X = 123 AND Y = 18 else
"111111111111" when X = 124 AND Y = 18 else
"111111111111" when X = 125 AND Y = 18 else
"111111111111" when X = 126 AND Y = 18 else
"111111111111" when X = 127 AND Y = 18 else
"111111111111" when X = 128 AND Y = 18 else
"111111111111" when X = 129 AND Y = 18 else
"111111111111" when X = 130 AND Y = 18 else
"111111111111" when X = 131 AND Y = 18 else
"111111111111" when X = 132 AND Y = 18 else
"111111111111" when X = 133 AND Y = 18 else
"111111111111" when X = 134 AND Y = 18 else
"111111111111" when X = 135 AND Y = 18 else
"111111111111" when X = 136 AND Y = 18 else
"111111111111" when X = 137 AND Y = 18 else
"111111111111" when X = 138 AND Y = 18 else
"111111111111" when X = 139 AND Y = 18 else
"111111111111" when X = 140 AND Y = 18 else
"111111111111" when X = 141 AND Y = 18 else
"111111111111" when X = 142 AND Y = 18 else
"111111111111" when X = 143 AND Y = 18 else
"111111111111" when X = 144 AND Y = 18 else
"111111111111" when X = 145 AND Y = 18 else
"111111111111" when X = 146 AND Y = 18 else
"111111111111" when X = 147 AND Y = 18 else
"111111111111" when X = 148 AND Y = 18 else
"111111111111" when X = 149 AND Y = 18 else
"111111111111" when X = 150 AND Y = 18 else
"111111111111" when X = 151 AND Y = 18 else
"111111111111" when X = 152 AND Y = 18 else
"111111111111" when X = 153 AND Y = 18 else
"111111111111" when X = 154 AND Y = 18 else
"000000000000" when X = 155 AND Y = 18 else
"000000000000" when X = 156 AND Y = 18 else
"000000000000" when X = 157 AND Y = 18 else
"000000000000" when X = 158 AND Y = 18 else
"000000000000" when X = 159 AND Y = 18 else
"000000000000" when X = 160 AND Y = 18 else
"000000000000" when X = 161 AND Y = 18 else
"000000000000" when X = 162 AND Y = 18 else
"000000000000" when X = 163 AND Y = 18 else
"000000000000" when X = 164 AND Y = 18 else
"000000000000" when X = 165 AND Y = 18 else
"000000000000" when X = 166 AND Y = 18 else
"000000000000" when X = 167 AND Y = 18 else
"000000000000" when X = 168 AND Y = 18 else
"000000000000" when X = 169 AND Y = 18 else
"000000000000" when X = 170 AND Y = 18 else
"000000000000" when X = 171 AND Y = 18 else
"000000000000" when X = 172 AND Y = 18 else
"000000000000" when X = 173 AND Y = 18 else
"000000000000" when X = 174 AND Y = 18 else
"000000000000" when X = 175 AND Y = 18 else
"000000000000" when X = 176 AND Y = 18 else
"000000000000" when X = 177 AND Y = 18 else
"000000000000" when X = 178 AND Y = 18 else
"000000000000" when X = 179 AND Y = 18 else
"000000000000" when X = 180 AND Y = 18 else
"000000000000" when X = 181 AND Y = 18 else
"000000000000" when X = 182 AND Y = 18 else
"000000000000" when X = 183 AND Y = 18 else
"000000000000" when X = 184 AND Y = 18 else
"000000000000" when X = 185 AND Y = 18 else
"000000000000" when X = 186 AND Y = 18 else
"000000000000" when X = 187 AND Y = 18 else
"000000000000" when X = 188 AND Y = 18 else
"000000000000" when X = 189 AND Y = 18 else
"000000000000" when X = 190 AND Y = 18 else
"000000000000" when X = 191 AND Y = 18 else
"000000000000" when X = 192 AND Y = 18 else
"000000000000" when X = 193 AND Y = 18 else
"000000000000" when X = 194 AND Y = 18 else
"000000000000" when X = 195 AND Y = 18 else
"000000000000" when X = 196 AND Y = 18 else
"000000000000" when X = 197 AND Y = 18 else
"000000000000" when X = 198 AND Y = 18 else
"000000000000" when X = 199 AND Y = 18 else
"000000000000" when X = 200 AND Y = 18 else
"000000000000" when X = 201 AND Y = 18 else
"000000000000" when X = 202 AND Y = 18 else
"000000000000" when X = 203 AND Y = 18 else
"000000000000" when X = 204 AND Y = 18 else
"000000000000" when X = 205 AND Y = 18 else
"000000000000" when X = 206 AND Y = 18 else
"000000000000" when X = 207 AND Y = 18 else
"000000000000" when X = 208 AND Y = 18 else
"000000000000" when X = 209 AND Y = 18 else
"000000000000" when X = 210 AND Y = 18 else
"000000000000" when X = 211 AND Y = 18 else
"000000000000" when X = 212 AND Y = 18 else
"000000000000" when X = 213 AND Y = 18 else
"000000000000" when X = 214 AND Y = 18 else
"000000000000" when X = 215 AND Y = 18 else
"000000000000" when X = 216 AND Y = 18 else
"000000000000" when X = 217 AND Y = 18 else
"000000000000" when X = 218 AND Y = 18 else
"000000000000" when X = 219 AND Y = 18 else
"000000000000" when X = 220 AND Y = 18 else
"000000000000" when X = 221 AND Y = 18 else
"000000000000" when X = 222 AND Y = 18 else
"000000000000" when X = 223 AND Y = 18 else
"000000000000" when X = 224 AND Y = 18 else
"000000000000" when X = 225 AND Y = 18 else
"000000000000" when X = 226 AND Y = 18 else
"000000000000" when X = 227 AND Y = 18 else
"000000000000" when X = 228 AND Y = 18 else
"000000000000" when X = 229 AND Y = 18 else
"000000000000" when X = 230 AND Y = 18 else
"000000000000" when X = 231 AND Y = 18 else
"000000000000" when X = 232 AND Y = 18 else
"000000000000" when X = 233 AND Y = 18 else
"000000000000" when X = 234 AND Y = 18 else
"000000000000" when X = 235 AND Y = 18 else
"000000000000" when X = 236 AND Y = 18 else
"000000000000" when X = 237 AND Y = 18 else
"000000000000" when X = 238 AND Y = 18 else
"000000000000" when X = 239 AND Y = 18 else
"000000000000" when X = 240 AND Y = 18 else
"000000000000" when X = 241 AND Y = 18 else
"000000000000" when X = 242 AND Y = 18 else
"000000000000" when X = 243 AND Y = 18 else
"000000000000" when X = 244 AND Y = 18 else
"000000000000" when X = 245 AND Y = 18 else
"000000000000" when X = 246 AND Y = 18 else
"000000000000" when X = 247 AND Y = 18 else
"000000000000" when X = 248 AND Y = 18 else
"000000000000" when X = 249 AND Y = 18 else
"000000000000" when X = 250 AND Y = 18 else
"000000000000" when X = 251 AND Y = 18 else
"000000000000" when X = 252 AND Y = 18 else
"000000000000" when X = 253 AND Y = 18 else
"000000000000" when X = 254 AND Y = 18 else
"000000000000" when X = 255 AND Y = 18 else
"000000000000" when X = 256 AND Y = 18 else
"000000000000" when X = 257 AND Y = 18 else
"000000000000" when X = 258 AND Y = 18 else
"000000000000" when X = 259 AND Y = 18 else
"000000000000" when X = 260 AND Y = 18 else
"000000000000" when X = 261 AND Y = 18 else
"000000000000" when X = 262 AND Y = 18 else
"000000000000" when X = 263 AND Y = 18 else
"000000000000" when X = 264 AND Y = 18 else
"000000000000" when X = 265 AND Y = 18 else
"000000000000" when X = 266 AND Y = 18 else
"000000000000" when X = 267 AND Y = 18 else
"000000000000" when X = 268 AND Y = 18 else
"000000000000" when X = 269 AND Y = 18 else
"000000000000" when X = 270 AND Y = 18 else
"000000000000" when X = 271 AND Y = 18 else
"000000000000" when X = 272 AND Y = 18 else
"000000000000" when X = 273 AND Y = 18 else
"000000000000" when X = 274 AND Y = 18 else
"000000000000" when X = 275 AND Y = 18 else
"000000000000" when X = 276 AND Y = 18 else
"000000000000" when X = 277 AND Y = 18 else
"000000000000" when X = 278 AND Y = 18 else
"000000000000" when X = 279 AND Y = 18 else
"000000000000" when X = 280 AND Y = 18 else
"000000000000" when X = 281 AND Y = 18 else
"000000000000" when X = 282 AND Y = 18 else
"000000000000" when X = 283 AND Y = 18 else
"000000000000" when X = 284 AND Y = 18 else
"000000000000" when X = 285 AND Y = 18 else
"000000000000" when X = 286 AND Y = 18 else
"000000000000" when X = 287 AND Y = 18 else
"000000000000" when X = 288 AND Y = 18 else
"000000000000" when X = 289 AND Y = 18 else
"000000000000" when X = 290 AND Y = 18 else
"000000000000" when X = 291 AND Y = 18 else
"000000000000" when X = 292 AND Y = 18 else
"000000000000" when X = 293 AND Y = 18 else
"000000000000" when X = 294 AND Y = 18 else
"000000000000" when X = 295 AND Y = 18 else
"000000000000" when X = 296 AND Y = 18 else
"000000000000" when X = 297 AND Y = 18 else
"000000000000" when X = 298 AND Y = 18 else
"000000000000" when X = 299 AND Y = 18 else
"000000000000" when X = 300 AND Y = 18 else
"000000000000" when X = 301 AND Y = 18 else
"000000000000" when X = 302 AND Y = 18 else
"000000000000" when X = 303 AND Y = 18 else
"000000000000" when X = 304 AND Y = 18 else
"000000000000" when X = 305 AND Y = 18 else
"000000000000" when X = 306 AND Y = 18 else
"000000000000" when X = 307 AND Y = 18 else
"000000000000" when X = 308 AND Y = 18 else
"000000000000" when X = 309 AND Y = 18 else
"000000000000" when X = 310 AND Y = 18 else
"000000000000" when X = 311 AND Y = 18 else
"000000000000" when X = 312 AND Y = 18 else
"000000000000" when X = 313 AND Y = 18 else
"000000000000" when X = 314 AND Y = 18 else
"000000000000" when X = 315 AND Y = 18 else
"000000000000" when X = 316 AND Y = 18 else
"000000000000" when X = 317 AND Y = 18 else
"000000000000" when X = 318 AND Y = 18 else
"000000000000" when X = 319 AND Y = 18 else
"000000000000" when X = 320 AND Y = 18 else
"000000000000" when X = 321 AND Y = 18 else
"000000000000" when X = 322 AND Y = 18 else
"000000000000" when X = 323 AND Y = 18 else
"000000000000" when X = 324 AND Y = 18 else
"000000000000" when X = 0 AND Y = 19 else
"000000000000" when X = 1 AND Y = 19 else
"000000000000" when X = 2 AND Y = 19 else
"000000000000" when X = 3 AND Y = 19 else
"000000000000" when X = 4 AND Y = 19 else
"000000000000" when X = 5 AND Y = 19 else
"000000000000" when X = 6 AND Y = 19 else
"000000000000" when X = 7 AND Y = 19 else
"000000000000" when X = 8 AND Y = 19 else
"000000000000" when X = 9 AND Y = 19 else
"000000000000" when X = 10 AND Y = 19 else
"000000000000" when X = 11 AND Y = 19 else
"000000000000" when X = 12 AND Y = 19 else
"000000000000" when X = 13 AND Y = 19 else
"000000000000" when X = 14 AND Y = 19 else
"000000000000" when X = 15 AND Y = 19 else
"000000000000" when X = 16 AND Y = 19 else
"000000000000" when X = 17 AND Y = 19 else
"000000000000" when X = 18 AND Y = 19 else
"000000000000" when X = 19 AND Y = 19 else
"000000000000" when X = 20 AND Y = 19 else
"000000000000" when X = 21 AND Y = 19 else
"000000000000" when X = 22 AND Y = 19 else
"000000000000" when X = 23 AND Y = 19 else
"000000000000" when X = 24 AND Y = 19 else
"000000000000" when X = 25 AND Y = 19 else
"000000000000" when X = 26 AND Y = 19 else
"000000000000" when X = 27 AND Y = 19 else
"000000000000" when X = 28 AND Y = 19 else
"000000000000" when X = 29 AND Y = 19 else
"000000000000" when X = 30 AND Y = 19 else
"000000000000" when X = 31 AND Y = 19 else
"000000000000" when X = 32 AND Y = 19 else
"000000000000" when X = 33 AND Y = 19 else
"000000000000" when X = 34 AND Y = 19 else
"000000000000" when X = 35 AND Y = 19 else
"000000000000" when X = 36 AND Y = 19 else
"000000000000" when X = 37 AND Y = 19 else
"000000000000" when X = 38 AND Y = 19 else
"000000000000" when X = 39 AND Y = 19 else
"100010011101" when X = 40 AND Y = 19 else
"100010011101" when X = 41 AND Y = 19 else
"100010011101" when X = 42 AND Y = 19 else
"100010011101" when X = 43 AND Y = 19 else
"100010011101" when X = 44 AND Y = 19 else
"100010011101" when X = 45 AND Y = 19 else
"100010011101" when X = 46 AND Y = 19 else
"100010011101" when X = 47 AND Y = 19 else
"100010011101" when X = 48 AND Y = 19 else
"100010011101" when X = 49 AND Y = 19 else
"110111011111" when X = 50 AND Y = 19 else
"110111011111" when X = 51 AND Y = 19 else
"110111011111" when X = 52 AND Y = 19 else
"110111011111" when X = 53 AND Y = 19 else
"110111011111" when X = 54 AND Y = 19 else
"110111011111" when X = 55 AND Y = 19 else
"110111011111" when X = 56 AND Y = 19 else
"110111011111" when X = 57 AND Y = 19 else
"110111011111" when X = 58 AND Y = 19 else
"110111011111" when X = 59 AND Y = 19 else
"110111011111" when X = 60 AND Y = 19 else
"110111011111" when X = 61 AND Y = 19 else
"110111011111" when X = 62 AND Y = 19 else
"110111011111" when X = 63 AND Y = 19 else
"110111011111" when X = 64 AND Y = 19 else
"111111111111" when X = 65 AND Y = 19 else
"111111111111" when X = 66 AND Y = 19 else
"111111111111" when X = 67 AND Y = 19 else
"111111111111" when X = 68 AND Y = 19 else
"111111111111" when X = 69 AND Y = 19 else
"111111111111" when X = 70 AND Y = 19 else
"111111111111" when X = 71 AND Y = 19 else
"111111111111" when X = 72 AND Y = 19 else
"111111111111" when X = 73 AND Y = 19 else
"111111111111" when X = 74 AND Y = 19 else
"111111111111" when X = 75 AND Y = 19 else
"111111111111" when X = 76 AND Y = 19 else
"111111111111" when X = 77 AND Y = 19 else
"111111111111" when X = 78 AND Y = 19 else
"111111111111" when X = 79 AND Y = 19 else
"111111111111" when X = 80 AND Y = 19 else
"111111111111" when X = 81 AND Y = 19 else
"111111111111" when X = 82 AND Y = 19 else
"111111111111" when X = 83 AND Y = 19 else
"111111111111" when X = 84 AND Y = 19 else
"111111111111" when X = 85 AND Y = 19 else
"111111111111" when X = 86 AND Y = 19 else
"111111111111" when X = 87 AND Y = 19 else
"111111111111" when X = 88 AND Y = 19 else
"111111111111" when X = 89 AND Y = 19 else
"111111111111" when X = 90 AND Y = 19 else
"111111111111" when X = 91 AND Y = 19 else
"111111111111" when X = 92 AND Y = 19 else
"111111111111" when X = 93 AND Y = 19 else
"111111111111" when X = 94 AND Y = 19 else
"111111111111" when X = 95 AND Y = 19 else
"111111111111" when X = 96 AND Y = 19 else
"111111111111" when X = 97 AND Y = 19 else
"111111111111" when X = 98 AND Y = 19 else
"111111111111" when X = 99 AND Y = 19 else
"111111111111" when X = 100 AND Y = 19 else
"111111111111" when X = 101 AND Y = 19 else
"111111111111" when X = 102 AND Y = 19 else
"111111111111" when X = 103 AND Y = 19 else
"111111111111" when X = 104 AND Y = 19 else
"111111111111" when X = 105 AND Y = 19 else
"111111111111" when X = 106 AND Y = 19 else
"111111111111" when X = 107 AND Y = 19 else
"111111111111" when X = 108 AND Y = 19 else
"111111111111" when X = 109 AND Y = 19 else
"111111111111" when X = 110 AND Y = 19 else
"111111111111" when X = 111 AND Y = 19 else
"111111111111" when X = 112 AND Y = 19 else
"111111111111" when X = 113 AND Y = 19 else
"111111111111" when X = 114 AND Y = 19 else
"111111111111" when X = 115 AND Y = 19 else
"111111111111" when X = 116 AND Y = 19 else
"111111111111" when X = 117 AND Y = 19 else
"111111111111" when X = 118 AND Y = 19 else
"111111111111" when X = 119 AND Y = 19 else
"111111111111" when X = 120 AND Y = 19 else
"111111111111" when X = 121 AND Y = 19 else
"111111111111" when X = 122 AND Y = 19 else
"111111111111" when X = 123 AND Y = 19 else
"111111111111" when X = 124 AND Y = 19 else
"111111111111" when X = 125 AND Y = 19 else
"111111111111" when X = 126 AND Y = 19 else
"111111111111" when X = 127 AND Y = 19 else
"111111111111" when X = 128 AND Y = 19 else
"111111111111" when X = 129 AND Y = 19 else
"111111111111" when X = 130 AND Y = 19 else
"111111111111" when X = 131 AND Y = 19 else
"111111111111" when X = 132 AND Y = 19 else
"111111111111" when X = 133 AND Y = 19 else
"111111111111" when X = 134 AND Y = 19 else
"111111111111" when X = 135 AND Y = 19 else
"111111111111" when X = 136 AND Y = 19 else
"111111111111" when X = 137 AND Y = 19 else
"111111111111" when X = 138 AND Y = 19 else
"111111111111" when X = 139 AND Y = 19 else
"111111111111" when X = 140 AND Y = 19 else
"111111111111" when X = 141 AND Y = 19 else
"111111111111" when X = 142 AND Y = 19 else
"111111111111" when X = 143 AND Y = 19 else
"111111111111" when X = 144 AND Y = 19 else
"111111111111" when X = 145 AND Y = 19 else
"111111111111" when X = 146 AND Y = 19 else
"111111111111" when X = 147 AND Y = 19 else
"111111111111" when X = 148 AND Y = 19 else
"111111111111" when X = 149 AND Y = 19 else
"111111111111" when X = 150 AND Y = 19 else
"111111111111" when X = 151 AND Y = 19 else
"111111111111" when X = 152 AND Y = 19 else
"111111111111" when X = 153 AND Y = 19 else
"111111111111" when X = 154 AND Y = 19 else
"000000000000" when X = 155 AND Y = 19 else
"000000000000" when X = 156 AND Y = 19 else
"000000000000" when X = 157 AND Y = 19 else
"000000000000" when X = 158 AND Y = 19 else
"000000000000" when X = 159 AND Y = 19 else
"000000000000" when X = 160 AND Y = 19 else
"000000000000" when X = 161 AND Y = 19 else
"000000000000" when X = 162 AND Y = 19 else
"000000000000" when X = 163 AND Y = 19 else
"000000000000" when X = 164 AND Y = 19 else
"000000000000" when X = 165 AND Y = 19 else
"000000000000" when X = 166 AND Y = 19 else
"000000000000" when X = 167 AND Y = 19 else
"000000000000" when X = 168 AND Y = 19 else
"000000000000" when X = 169 AND Y = 19 else
"000000000000" when X = 170 AND Y = 19 else
"000000000000" when X = 171 AND Y = 19 else
"000000000000" when X = 172 AND Y = 19 else
"000000000000" when X = 173 AND Y = 19 else
"000000000000" when X = 174 AND Y = 19 else
"000000000000" when X = 175 AND Y = 19 else
"000000000000" when X = 176 AND Y = 19 else
"000000000000" when X = 177 AND Y = 19 else
"000000000000" when X = 178 AND Y = 19 else
"000000000000" when X = 179 AND Y = 19 else
"000000000000" when X = 180 AND Y = 19 else
"000000000000" when X = 181 AND Y = 19 else
"000000000000" when X = 182 AND Y = 19 else
"000000000000" when X = 183 AND Y = 19 else
"000000000000" when X = 184 AND Y = 19 else
"000000000000" when X = 185 AND Y = 19 else
"000000000000" when X = 186 AND Y = 19 else
"000000000000" when X = 187 AND Y = 19 else
"000000000000" when X = 188 AND Y = 19 else
"000000000000" when X = 189 AND Y = 19 else
"000000000000" when X = 190 AND Y = 19 else
"000000000000" when X = 191 AND Y = 19 else
"000000000000" when X = 192 AND Y = 19 else
"000000000000" when X = 193 AND Y = 19 else
"000000000000" when X = 194 AND Y = 19 else
"000000000000" when X = 195 AND Y = 19 else
"000000000000" when X = 196 AND Y = 19 else
"000000000000" when X = 197 AND Y = 19 else
"000000000000" when X = 198 AND Y = 19 else
"000000000000" when X = 199 AND Y = 19 else
"000000000000" when X = 200 AND Y = 19 else
"000000000000" when X = 201 AND Y = 19 else
"000000000000" when X = 202 AND Y = 19 else
"000000000000" when X = 203 AND Y = 19 else
"000000000000" when X = 204 AND Y = 19 else
"000000000000" when X = 205 AND Y = 19 else
"000000000000" when X = 206 AND Y = 19 else
"000000000000" when X = 207 AND Y = 19 else
"000000000000" when X = 208 AND Y = 19 else
"000000000000" when X = 209 AND Y = 19 else
"000000000000" when X = 210 AND Y = 19 else
"000000000000" when X = 211 AND Y = 19 else
"000000000000" when X = 212 AND Y = 19 else
"000000000000" when X = 213 AND Y = 19 else
"000000000000" when X = 214 AND Y = 19 else
"000000000000" when X = 215 AND Y = 19 else
"000000000000" when X = 216 AND Y = 19 else
"000000000000" when X = 217 AND Y = 19 else
"000000000000" when X = 218 AND Y = 19 else
"000000000000" when X = 219 AND Y = 19 else
"000000000000" when X = 220 AND Y = 19 else
"000000000000" when X = 221 AND Y = 19 else
"000000000000" when X = 222 AND Y = 19 else
"000000000000" when X = 223 AND Y = 19 else
"000000000000" when X = 224 AND Y = 19 else
"000000000000" when X = 225 AND Y = 19 else
"000000000000" when X = 226 AND Y = 19 else
"000000000000" when X = 227 AND Y = 19 else
"000000000000" when X = 228 AND Y = 19 else
"000000000000" when X = 229 AND Y = 19 else
"000000000000" when X = 230 AND Y = 19 else
"000000000000" when X = 231 AND Y = 19 else
"000000000000" when X = 232 AND Y = 19 else
"000000000000" when X = 233 AND Y = 19 else
"000000000000" when X = 234 AND Y = 19 else
"000000000000" when X = 235 AND Y = 19 else
"000000000000" when X = 236 AND Y = 19 else
"000000000000" when X = 237 AND Y = 19 else
"000000000000" when X = 238 AND Y = 19 else
"000000000000" when X = 239 AND Y = 19 else
"000000000000" when X = 240 AND Y = 19 else
"000000000000" when X = 241 AND Y = 19 else
"000000000000" when X = 242 AND Y = 19 else
"000000000000" when X = 243 AND Y = 19 else
"000000000000" when X = 244 AND Y = 19 else
"000000000000" when X = 245 AND Y = 19 else
"000000000000" when X = 246 AND Y = 19 else
"000000000000" when X = 247 AND Y = 19 else
"000000000000" when X = 248 AND Y = 19 else
"000000000000" when X = 249 AND Y = 19 else
"000000000000" when X = 250 AND Y = 19 else
"000000000000" when X = 251 AND Y = 19 else
"000000000000" when X = 252 AND Y = 19 else
"000000000000" when X = 253 AND Y = 19 else
"000000000000" when X = 254 AND Y = 19 else
"000000000000" when X = 255 AND Y = 19 else
"000000000000" when X = 256 AND Y = 19 else
"000000000000" when X = 257 AND Y = 19 else
"000000000000" when X = 258 AND Y = 19 else
"000000000000" when X = 259 AND Y = 19 else
"000000000000" when X = 260 AND Y = 19 else
"000000000000" when X = 261 AND Y = 19 else
"000000000000" when X = 262 AND Y = 19 else
"000000000000" when X = 263 AND Y = 19 else
"000000000000" when X = 264 AND Y = 19 else
"000000000000" when X = 265 AND Y = 19 else
"000000000000" when X = 266 AND Y = 19 else
"000000000000" when X = 267 AND Y = 19 else
"000000000000" when X = 268 AND Y = 19 else
"000000000000" when X = 269 AND Y = 19 else
"000000000000" when X = 270 AND Y = 19 else
"000000000000" when X = 271 AND Y = 19 else
"000000000000" when X = 272 AND Y = 19 else
"000000000000" when X = 273 AND Y = 19 else
"000000000000" when X = 274 AND Y = 19 else
"000000000000" when X = 275 AND Y = 19 else
"000000000000" when X = 276 AND Y = 19 else
"000000000000" when X = 277 AND Y = 19 else
"000000000000" when X = 278 AND Y = 19 else
"000000000000" when X = 279 AND Y = 19 else
"000000000000" when X = 280 AND Y = 19 else
"000000000000" when X = 281 AND Y = 19 else
"000000000000" when X = 282 AND Y = 19 else
"000000000000" when X = 283 AND Y = 19 else
"000000000000" when X = 284 AND Y = 19 else
"000000000000" when X = 285 AND Y = 19 else
"000000000000" when X = 286 AND Y = 19 else
"000000000000" when X = 287 AND Y = 19 else
"000000000000" when X = 288 AND Y = 19 else
"000000000000" when X = 289 AND Y = 19 else
"000000000000" when X = 290 AND Y = 19 else
"000000000000" when X = 291 AND Y = 19 else
"000000000000" when X = 292 AND Y = 19 else
"000000000000" when X = 293 AND Y = 19 else
"000000000000" when X = 294 AND Y = 19 else
"000000000000" when X = 295 AND Y = 19 else
"000000000000" when X = 296 AND Y = 19 else
"000000000000" when X = 297 AND Y = 19 else
"000000000000" when X = 298 AND Y = 19 else
"000000000000" when X = 299 AND Y = 19 else
"000000000000" when X = 300 AND Y = 19 else
"000000000000" when X = 301 AND Y = 19 else
"000000000000" when X = 302 AND Y = 19 else
"000000000000" when X = 303 AND Y = 19 else
"000000000000" when X = 304 AND Y = 19 else
"000000000000" when X = 305 AND Y = 19 else
"000000000000" when X = 306 AND Y = 19 else
"000000000000" when X = 307 AND Y = 19 else
"000000000000" when X = 308 AND Y = 19 else
"000000000000" when X = 309 AND Y = 19 else
"000000000000" when X = 310 AND Y = 19 else
"000000000000" when X = 311 AND Y = 19 else
"000000000000" when X = 312 AND Y = 19 else
"000000000000" when X = 313 AND Y = 19 else
"000000000000" when X = 314 AND Y = 19 else
"000000000000" when X = 315 AND Y = 19 else
"000000000000" when X = 316 AND Y = 19 else
"000000000000" when X = 317 AND Y = 19 else
"000000000000" when X = 318 AND Y = 19 else
"000000000000" when X = 319 AND Y = 19 else
"000000000000" when X = 320 AND Y = 19 else
"000000000000" when X = 321 AND Y = 19 else
"000000000000" when X = 322 AND Y = 19 else
"000000000000" when X = 323 AND Y = 19 else
"000000000000" when X = 324 AND Y = 19 else
"000000000000" when X = 0 AND Y = 20 else
"000000000000" when X = 1 AND Y = 20 else
"000000000000" when X = 2 AND Y = 20 else
"000000000000" when X = 3 AND Y = 20 else
"000000000000" when X = 4 AND Y = 20 else
"000000000000" when X = 5 AND Y = 20 else
"000000000000" when X = 6 AND Y = 20 else
"000000000000" when X = 7 AND Y = 20 else
"000000000000" when X = 8 AND Y = 20 else
"000000000000" when X = 9 AND Y = 20 else
"000000000000" when X = 10 AND Y = 20 else
"000000000000" when X = 11 AND Y = 20 else
"000000000000" when X = 12 AND Y = 20 else
"000000000000" when X = 13 AND Y = 20 else
"000000000000" when X = 14 AND Y = 20 else
"000000000000" when X = 15 AND Y = 20 else
"000000000000" when X = 16 AND Y = 20 else
"000000000000" when X = 17 AND Y = 20 else
"000000000000" when X = 18 AND Y = 20 else
"000000000000" when X = 19 AND Y = 20 else
"000000000000" when X = 20 AND Y = 20 else
"000000000000" when X = 21 AND Y = 20 else
"000000000000" when X = 22 AND Y = 20 else
"000000000000" when X = 23 AND Y = 20 else
"000000000000" when X = 24 AND Y = 20 else
"000000000000" when X = 25 AND Y = 20 else
"000000000000" when X = 26 AND Y = 20 else
"000000000000" when X = 27 AND Y = 20 else
"000000000000" when X = 28 AND Y = 20 else
"000000000000" when X = 29 AND Y = 20 else
"000000000000" when X = 30 AND Y = 20 else
"000000000000" when X = 31 AND Y = 20 else
"000000000000" when X = 32 AND Y = 20 else
"000000000000" when X = 33 AND Y = 20 else
"000000000000" when X = 34 AND Y = 20 else
"000000000000" when X = 35 AND Y = 20 else
"000000000000" when X = 36 AND Y = 20 else
"000000000000" when X = 37 AND Y = 20 else
"000000000000" when X = 38 AND Y = 20 else
"000000000000" when X = 39 AND Y = 20 else
"100010011101" when X = 40 AND Y = 20 else
"100010011101" when X = 41 AND Y = 20 else
"100010011101" when X = 42 AND Y = 20 else
"100010011101" when X = 43 AND Y = 20 else
"100010011101" when X = 44 AND Y = 20 else
"100010011101" when X = 45 AND Y = 20 else
"100010011101" when X = 46 AND Y = 20 else
"100010011101" when X = 47 AND Y = 20 else
"100010011101" when X = 48 AND Y = 20 else
"100010011101" when X = 49 AND Y = 20 else
"110111011111" when X = 50 AND Y = 20 else
"110111011111" when X = 51 AND Y = 20 else
"110111011111" when X = 52 AND Y = 20 else
"110111011111" when X = 53 AND Y = 20 else
"110111011111" when X = 54 AND Y = 20 else
"110111011111" when X = 55 AND Y = 20 else
"110111011111" when X = 56 AND Y = 20 else
"110111011111" when X = 57 AND Y = 20 else
"110111011111" when X = 58 AND Y = 20 else
"110111011111" when X = 59 AND Y = 20 else
"111111111111" when X = 60 AND Y = 20 else
"111111111111" when X = 61 AND Y = 20 else
"111111111111" when X = 62 AND Y = 20 else
"111111111111" when X = 63 AND Y = 20 else
"111111111111" when X = 64 AND Y = 20 else
"111111111111" when X = 65 AND Y = 20 else
"111111111111" when X = 66 AND Y = 20 else
"111111111111" when X = 67 AND Y = 20 else
"111111111111" when X = 68 AND Y = 20 else
"111111111111" when X = 69 AND Y = 20 else
"111111111111" when X = 70 AND Y = 20 else
"111111111111" when X = 71 AND Y = 20 else
"111111111111" when X = 72 AND Y = 20 else
"111111111111" when X = 73 AND Y = 20 else
"111111111111" when X = 74 AND Y = 20 else
"111111111111" when X = 75 AND Y = 20 else
"111111111111" when X = 76 AND Y = 20 else
"111111111111" when X = 77 AND Y = 20 else
"111111111111" when X = 78 AND Y = 20 else
"111111111111" when X = 79 AND Y = 20 else
"111111111111" when X = 80 AND Y = 20 else
"111111111111" when X = 81 AND Y = 20 else
"111111111111" when X = 82 AND Y = 20 else
"111111111111" when X = 83 AND Y = 20 else
"111111111111" when X = 84 AND Y = 20 else
"111111111111" when X = 85 AND Y = 20 else
"111111111111" when X = 86 AND Y = 20 else
"111111111111" when X = 87 AND Y = 20 else
"111111111111" when X = 88 AND Y = 20 else
"111111111111" when X = 89 AND Y = 20 else
"111111111111" when X = 90 AND Y = 20 else
"111111111111" when X = 91 AND Y = 20 else
"111111111111" when X = 92 AND Y = 20 else
"111111111111" when X = 93 AND Y = 20 else
"111111111111" when X = 94 AND Y = 20 else
"111111111111" when X = 95 AND Y = 20 else
"111111111111" when X = 96 AND Y = 20 else
"111111111111" when X = 97 AND Y = 20 else
"111111111111" when X = 98 AND Y = 20 else
"111111111111" when X = 99 AND Y = 20 else
"111111111111" when X = 100 AND Y = 20 else
"111111111111" when X = 101 AND Y = 20 else
"111111111111" when X = 102 AND Y = 20 else
"111111111111" when X = 103 AND Y = 20 else
"111111111111" when X = 104 AND Y = 20 else
"111111111111" when X = 105 AND Y = 20 else
"111111111111" when X = 106 AND Y = 20 else
"111111111111" when X = 107 AND Y = 20 else
"111111111111" when X = 108 AND Y = 20 else
"111111111111" when X = 109 AND Y = 20 else
"111111111111" when X = 110 AND Y = 20 else
"111111111111" when X = 111 AND Y = 20 else
"111111111111" when X = 112 AND Y = 20 else
"111111111111" when X = 113 AND Y = 20 else
"111111111111" when X = 114 AND Y = 20 else
"111111111111" when X = 115 AND Y = 20 else
"111111111111" when X = 116 AND Y = 20 else
"111111111111" when X = 117 AND Y = 20 else
"111111111111" when X = 118 AND Y = 20 else
"111111111111" when X = 119 AND Y = 20 else
"111111111111" when X = 120 AND Y = 20 else
"111111111111" when X = 121 AND Y = 20 else
"111111111111" when X = 122 AND Y = 20 else
"111111111111" when X = 123 AND Y = 20 else
"111111111111" when X = 124 AND Y = 20 else
"111111111111" when X = 125 AND Y = 20 else
"111111111111" when X = 126 AND Y = 20 else
"111111111111" when X = 127 AND Y = 20 else
"111111111111" when X = 128 AND Y = 20 else
"111111111111" when X = 129 AND Y = 20 else
"111111111111" when X = 130 AND Y = 20 else
"111111111111" when X = 131 AND Y = 20 else
"111111111111" when X = 132 AND Y = 20 else
"111111111111" when X = 133 AND Y = 20 else
"111111111111" when X = 134 AND Y = 20 else
"111111111111" when X = 135 AND Y = 20 else
"111111111111" when X = 136 AND Y = 20 else
"111111111111" when X = 137 AND Y = 20 else
"111111111111" when X = 138 AND Y = 20 else
"111111111111" when X = 139 AND Y = 20 else
"111111111111" when X = 140 AND Y = 20 else
"111111111111" when X = 141 AND Y = 20 else
"111111111111" when X = 142 AND Y = 20 else
"111111111111" when X = 143 AND Y = 20 else
"111111111111" when X = 144 AND Y = 20 else
"111111111111" when X = 145 AND Y = 20 else
"111111111111" when X = 146 AND Y = 20 else
"111111111111" when X = 147 AND Y = 20 else
"111111111111" when X = 148 AND Y = 20 else
"111111111111" when X = 149 AND Y = 20 else
"111111111111" when X = 150 AND Y = 20 else
"111111111111" when X = 151 AND Y = 20 else
"111111111111" when X = 152 AND Y = 20 else
"111111111111" when X = 153 AND Y = 20 else
"111111111111" when X = 154 AND Y = 20 else
"000000000000" when X = 155 AND Y = 20 else
"000000000000" when X = 156 AND Y = 20 else
"000000000000" when X = 157 AND Y = 20 else
"000000000000" when X = 158 AND Y = 20 else
"000000000000" when X = 159 AND Y = 20 else
"000000000000" when X = 160 AND Y = 20 else
"000000000000" when X = 161 AND Y = 20 else
"000000000000" when X = 162 AND Y = 20 else
"000000000000" when X = 163 AND Y = 20 else
"000000000000" when X = 164 AND Y = 20 else
"000000000000" when X = 165 AND Y = 20 else
"000000000000" when X = 166 AND Y = 20 else
"000000000000" when X = 167 AND Y = 20 else
"000000000000" when X = 168 AND Y = 20 else
"000000000000" when X = 169 AND Y = 20 else
"000000000000" when X = 170 AND Y = 20 else
"000000000000" when X = 171 AND Y = 20 else
"000000000000" when X = 172 AND Y = 20 else
"000000000000" when X = 173 AND Y = 20 else
"000000000000" when X = 174 AND Y = 20 else
"000000000000" when X = 175 AND Y = 20 else
"000000000000" when X = 176 AND Y = 20 else
"000000000000" when X = 177 AND Y = 20 else
"000000000000" when X = 178 AND Y = 20 else
"000000000000" when X = 179 AND Y = 20 else
"000000000000" when X = 180 AND Y = 20 else
"000000000000" when X = 181 AND Y = 20 else
"000000000000" when X = 182 AND Y = 20 else
"000000000000" when X = 183 AND Y = 20 else
"000000000000" when X = 184 AND Y = 20 else
"000000000000" when X = 185 AND Y = 20 else
"000000000000" when X = 186 AND Y = 20 else
"000000000000" when X = 187 AND Y = 20 else
"000000000000" when X = 188 AND Y = 20 else
"000000000000" when X = 189 AND Y = 20 else
"000000000000" when X = 190 AND Y = 20 else
"000000000000" when X = 191 AND Y = 20 else
"000000000000" when X = 192 AND Y = 20 else
"000000000000" when X = 193 AND Y = 20 else
"000000000000" when X = 194 AND Y = 20 else
"000000000000" when X = 195 AND Y = 20 else
"000000000000" when X = 196 AND Y = 20 else
"000000000000" when X = 197 AND Y = 20 else
"000000000000" when X = 198 AND Y = 20 else
"000000000000" when X = 199 AND Y = 20 else
"000000000000" when X = 200 AND Y = 20 else
"000000000000" when X = 201 AND Y = 20 else
"000000000000" when X = 202 AND Y = 20 else
"000000000000" when X = 203 AND Y = 20 else
"000000000000" when X = 204 AND Y = 20 else
"000000000000" when X = 205 AND Y = 20 else
"000000000000" when X = 206 AND Y = 20 else
"000000000000" when X = 207 AND Y = 20 else
"000000000000" when X = 208 AND Y = 20 else
"000000000000" when X = 209 AND Y = 20 else
"000000000000" when X = 210 AND Y = 20 else
"000000000000" when X = 211 AND Y = 20 else
"000000000000" when X = 212 AND Y = 20 else
"000000000000" when X = 213 AND Y = 20 else
"000000000000" when X = 214 AND Y = 20 else
"000000000000" when X = 215 AND Y = 20 else
"000000000000" when X = 216 AND Y = 20 else
"000000000000" when X = 217 AND Y = 20 else
"000000000000" when X = 218 AND Y = 20 else
"000000000000" when X = 219 AND Y = 20 else
"000000000000" when X = 220 AND Y = 20 else
"000000000000" when X = 221 AND Y = 20 else
"000000000000" when X = 222 AND Y = 20 else
"000000000000" when X = 223 AND Y = 20 else
"000000000000" when X = 224 AND Y = 20 else
"000000000000" when X = 225 AND Y = 20 else
"000000000000" when X = 226 AND Y = 20 else
"000000000000" when X = 227 AND Y = 20 else
"000000000000" when X = 228 AND Y = 20 else
"000000000000" when X = 229 AND Y = 20 else
"000000000000" when X = 230 AND Y = 20 else
"000000000000" when X = 231 AND Y = 20 else
"000000000000" when X = 232 AND Y = 20 else
"000000000000" when X = 233 AND Y = 20 else
"000000000000" when X = 234 AND Y = 20 else
"000000000000" when X = 235 AND Y = 20 else
"000000000000" when X = 236 AND Y = 20 else
"000000000000" when X = 237 AND Y = 20 else
"000000000000" when X = 238 AND Y = 20 else
"000000000000" when X = 239 AND Y = 20 else
"000000000000" when X = 240 AND Y = 20 else
"000000000000" when X = 241 AND Y = 20 else
"000000000000" when X = 242 AND Y = 20 else
"000000000000" when X = 243 AND Y = 20 else
"000000000000" when X = 244 AND Y = 20 else
"000000000000" when X = 245 AND Y = 20 else
"000000000000" when X = 246 AND Y = 20 else
"000000000000" when X = 247 AND Y = 20 else
"000000000000" when X = 248 AND Y = 20 else
"000000000000" when X = 249 AND Y = 20 else
"000000000000" when X = 250 AND Y = 20 else
"000000000000" when X = 251 AND Y = 20 else
"000000000000" when X = 252 AND Y = 20 else
"000000000000" when X = 253 AND Y = 20 else
"000000000000" when X = 254 AND Y = 20 else
"000000000000" when X = 255 AND Y = 20 else
"000000000000" when X = 256 AND Y = 20 else
"000000000000" when X = 257 AND Y = 20 else
"000000000000" when X = 258 AND Y = 20 else
"000000000000" when X = 259 AND Y = 20 else
"000000000000" when X = 260 AND Y = 20 else
"000000000000" when X = 261 AND Y = 20 else
"000000000000" when X = 262 AND Y = 20 else
"000000000000" when X = 263 AND Y = 20 else
"000000000000" when X = 264 AND Y = 20 else
"000000000000" when X = 265 AND Y = 20 else
"000000000000" when X = 266 AND Y = 20 else
"000000000000" when X = 267 AND Y = 20 else
"000000000000" when X = 268 AND Y = 20 else
"000000000000" when X = 269 AND Y = 20 else
"000000000000" when X = 270 AND Y = 20 else
"000000000000" when X = 271 AND Y = 20 else
"000000000000" when X = 272 AND Y = 20 else
"000000000000" when X = 273 AND Y = 20 else
"000000000000" when X = 274 AND Y = 20 else
"000000000000" when X = 275 AND Y = 20 else
"000000000000" when X = 276 AND Y = 20 else
"000000000000" when X = 277 AND Y = 20 else
"000000000000" when X = 278 AND Y = 20 else
"000000000000" when X = 279 AND Y = 20 else
"000000000000" when X = 280 AND Y = 20 else
"000000000000" when X = 281 AND Y = 20 else
"000000000000" when X = 282 AND Y = 20 else
"000000000000" when X = 283 AND Y = 20 else
"000000000000" when X = 284 AND Y = 20 else
"000000000000" when X = 285 AND Y = 20 else
"000000000000" when X = 286 AND Y = 20 else
"000000000000" when X = 287 AND Y = 20 else
"000000000000" when X = 288 AND Y = 20 else
"000000000000" when X = 289 AND Y = 20 else
"000000000000" when X = 290 AND Y = 20 else
"000000000000" when X = 291 AND Y = 20 else
"000000000000" when X = 292 AND Y = 20 else
"000000000000" when X = 293 AND Y = 20 else
"000000000000" when X = 294 AND Y = 20 else
"000000000000" when X = 295 AND Y = 20 else
"000000000000" when X = 296 AND Y = 20 else
"000000000000" when X = 297 AND Y = 20 else
"000000000000" when X = 298 AND Y = 20 else
"000000000000" when X = 299 AND Y = 20 else
"000000000000" when X = 300 AND Y = 20 else
"000000000000" when X = 301 AND Y = 20 else
"000000000000" when X = 302 AND Y = 20 else
"000000000000" when X = 303 AND Y = 20 else
"000000000000" when X = 304 AND Y = 20 else
"000000000000" when X = 305 AND Y = 20 else
"000000000000" when X = 306 AND Y = 20 else
"000000000000" when X = 307 AND Y = 20 else
"000000000000" when X = 308 AND Y = 20 else
"000000000000" when X = 309 AND Y = 20 else
"000000000000" when X = 310 AND Y = 20 else
"000000000000" when X = 311 AND Y = 20 else
"000000000000" when X = 312 AND Y = 20 else
"000000000000" when X = 313 AND Y = 20 else
"000000000000" when X = 314 AND Y = 20 else
"000000000000" when X = 315 AND Y = 20 else
"000000000000" when X = 316 AND Y = 20 else
"000000000000" when X = 317 AND Y = 20 else
"000000000000" when X = 318 AND Y = 20 else
"000000000000" when X = 319 AND Y = 20 else
"000000000000" when X = 320 AND Y = 20 else
"000000000000" when X = 321 AND Y = 20 else
"000000000000" when X = 322 AND Y = 20 else
"000000000000" when X = 323 AND Y = 20 else
"000000000000" when X = 324 AND Y = 20 else
"000000000000" when X = 0 AND Y = 21 else
"000000000000" when X = 1 AND Y = 21 else
"000000000000" when X = 2 AND Y = 21 else
"000000000000" when X = 3 AND Y = 21 else
"000000000000" when X = 4 AND Y = 21 else
"000000000000" when X = 5 AND Y = 21 else
"000000000000" when X = 6 AND Y = 21 else
"000000000000" when X = 7 AND Y = 21 else
"000000000000" when X = 8 AND Y = 21 else
"000000000000" when X = 9 AND Y = 21 else
"000000000000" when X = 10 AND Y = 21 else
"000000000000" when X = 11 AND Y = 21 else
"000000000000" when X = 12 AND Y = 21 else
"000000000000" when X = 13 AND Y = 21 else
"000000000000" when X = 14 AND Y = 21 else
"000000000000" when X = 15 AND Y = 21 else
"000000000000" when X = 16 AND Y = 21 else
"000000000000" when X = 17 AND Y = 21 else
"000000000000" when X = 18 AND Y = 21 else
"000000000000" when X = 19 AND Y = 21 else
"000000000000" when X = 20 AND Y = 21 else
"000000000000" when X = 21 AND Y = 21 else
"000000000000" when X = 22 AND Y = 21 else
"000000000000" when X = 23 AND Y = 21 else
"000000000000" when X = 24 AND Y = 21 else
"000000000000" when X = 25 AND Y = 21 else
"000000000000" when X = 26 AND Y = 21 else
"000000000000" when X = 27 AND Y = 21 else
"000000000000" when X = 28 AND Y = 21 else
"000000000000" when X = 29 AND Y = 21 else
"000000000000" when X = 30 AND Y = 21 else
"000000000000" when X = 31 AND Y = 21 else
"000000000000" when X = 32 AND Y = 21 else
"000000000000" when X = 33 AND Y = 21 else
"000000000000" when X = 34 AND Y = 21 else
"000000000000" when X = 35 AND Y = 21 else
"000000000000" when X = 36 AND Y = 21 else
"000000000000" when X = 37 AND Y = 21 else
"000000000000" when X = 38 AND Y = 21 else
"000000000000" when X = 39 AND Y = 21 else
"100010011101" when X = 40 AND Y = 21 else
"100010011101" when X = 41 AND Y = 21 else
"100010011101" when X = 42 AND Y = 21 else
"100010011101" when X = 43 AND Y = 21 else
"100010011101" when X = 44 AND Y = 21 else
"100010011101" when X = 45 AND Y = 21 else
"100010011101" when X = 46 AND Y = 21 else
"100010011101" when X = 47 AND Y = 21 else
"100010011101" when X = 48 AND Y = 21 else
"100010011101" when X = 49 AND Y = 21 else
"110111011111" when X = 50 AND Y = 21 else
"110111011111" when X = 51 AND Y = 21 else
"110111011111" when X = 52 AND Y = 21 else
"110111011111" when X = 53 AND Y = 21 else
"110111011111" when X = 54 AND Y = 21 else
"110111011111" when X = 55 AND Y = 21 else
"110111011111" when X = 56 AND Y = 21 else
"110111011111" when X = 57 AND Y = 21 else
"110111011111" when X = 58 AND Y = 21 else
"110111011111" when X = 59 AND Y = 21 else
"111111111111" when X = 60 AND Y = 21 else
"111111111111" when X = 61 AND Y = 21 else
"111111111111" when X = 62 AND Y = 21 else
"111111111111" when X = 63 AND Y = 21 else
"111111111111" when X = 64 AND Y = 21 else
"111111111111" when X = 65 AND Y = 21 else
"111111111111" when X = 66 AND Y = 21 else
"111111111111" when X = 67 AND Y = 21 else
"111111111111" when X = 68 AND Y = 21 else
"111111111111" when X = 69 AND Y = 21 else
"111111111111" when X = 70 AND Y = 21 else
"111111111111" when X = 71 AND Y = 21 else
"111111111111" when X = 72 AND Y = 21 else
"111111111111" when X = 73 AND Y = 21 else
"111111111111" when X = 74 AND Y = 21 else
"111111111111" when X = 75 AND Y = 21 else
"111111111111" when X = 76 AND Y = 21 else
"111111111111" when X = 77 AND Y = 21 else
"111111111111" when X = 78 AND Y = 21 else
"111111111111" when X = 79 AND Y = 21 else
"111111111111" when X = 80 AND Y = 21 else
"111111111111" when X = 81 AND Y = 21 else
"111111111111" when X = 82 AND Y = 21 else
"111111111111" when X = 83 AND Y = 21 else
"111111111111" when X = 84 AND Y = 21 else
"111111111111" when X = 85 AND Y = 21 else
"111111111111" when X = 86 AND Y = 21 else
"111111111111" when X = 87 AND Y = 21 else
"111111111111" when X = 88 AND Y = 21 else
"111111111111" when X = 89 AND Y = 21 else
"111111111111" when X = 90 AND Y = 21 else
"111111111111" when X = 91 AND Y = 21 else
"111111111111" when X = 92 AND Y = 21 else
"111111111111" when X = 93 AND Y = 21 else
"111111111111" when X = 94 AND Y = 21 else
"111111111111" when X = 95 AND Y = 21 else
"111111111111" when X = 96 AND Y = 21 else
"111111111111" when X = 97 AND Y = 21 else
"111111111111" when X = 98 AND Y = 21 else
"111111111111" when X = 99 AND Y = 21 else
"111111111111" when X = 100 AND Y = 21 else
"111111111111" when X = 101 AND Y = 21 else
"111111111111" when X = 102 AND Y = 21 else
"111111111111" when X = 103 AND Y = 21 else
"111111111111" when X = 104 AND Y = 21 else
"111111111111" when X = 105 AND Y = 21 else
"111111111111" when X = 106 AND Y = 21 else
"111111111111" when X = 107 AND Y = 21 else
"111111111111" when X = 108 AND Y = 21 else
"111111111111" when X = 109 AND Y = 21 else
"111111111111" when X = 110 AND Y = 21 else
"111111111111" when X = 111 AND Y = 21 else
"111111111111" when X = 112 AND Y = 21 else
"111111111111" when X = 113 AND Y = 21 else
"111111111111" when X = 114 AND Y = 21 else
"111111111111" when X = 115 AND Y = 21 else
"111111111111" when X = 116 AND Y = 21 else
"111111111111" when X = 117 AND Y = 21 else
"111111111111" when X = 118 AND Y = 21 else
"111111111111" when X = 119 AND Y = 21 else
"111111111111" when X = 120 AND Y = 21 else
"111111111111" when X = 121 AND Y = 21 else
"111111111111" when X = 122 AND Y = 21 else
"111111111111" when X = 123 AND Y = 21 else
"111111111111" when X = 124 AND Y = 21 else
"111111111111" when X = 125 AND Y = 21 else
"111111111111" when X = 126 AND Y = 21 else
"111111111111" when X = 127 AND Y = 21 else
"111111111111" when X = 128 AND Y = 21 else
"111111111111" when X = 129 AND Y = 21 else
"111111111111" when X = 130 AND Y = 21 else
"111111111111" when X = 131 AND Y = 21 else
"111111111111" when X = 132 AND Y = 21 else
"111111111111" when X = 133 AND Y = 21 else
"111111111111" when X = 134 AND Y = 21 else
"111111111111" when X = 135 AND Y = 21 else
"111111111111" when X = 136 AND Y = 21 else
"111111111111" when X = 137 AND Y = 21 else
"111111111111" when X = 138 AND Y = 21 else
"111111111111" when X = 139 AND Y = 21 else
"111111111111" when X = 140 AND Y = 21 else
"111111111111" when X = 141 AND Y = 21 else
"111111111111" when X = 142 AND Y = 21 else
"111111111111" when X = 143 AND Y = 21 else
"111111111111" when X = 144 AND Y = 21 else
"111111111111" when X = 145 AND Y = 21 else
"111111111111" when X = 146 AND Y = 21 else
"111111111111" when X = 147 AND Y = 21 else
"111111111111" when X = 148 AND Y = 21 else
"111111111111" when X = 149 AND Y = 21 else
"111111111111" when X = 150 AND Y = 21 else
"111111111111" when X = 151 AND Y = 21 else
"111111111111" when X = 152 AND Y = 21 else
"111111111111" when X = 153 AND Y = 21 else
"111111111111" when X = 154 AND Y = 21 else
"000000000000" when X = 155 AND Y = 21 else
"000000000000" when X = 156 AND Y = 21 else
"000000000000" when X = 157 AND Y = 21 else
"000000000000" when X = 158 AND Y = 21 else
"000000000000" when X = 159 AND Y = 21 else
"000000000000" when X = 160 AND Y = 21 else
"000000000000" when X = 161 AND Y = 21 else
"000000000000" when X = 162 AND Y = 21 else
"000000000000" when X = 163 AND Y = 21 else
"000000000000" when X = 164 AND Y = 21 else
"000000000000" when X = 165 AND Y = 21 else
"000000000000" when X = 166 AND Y = 21 else
"000000000000" when X = 167 AND Y = 21 else
"000000000000" when X = 168 AND Y = 21 else
"000000000000" when X = 169 AND Y = 21 else
"000000000000" when X = 170 AND Y = 21 else
"000000000000" when X = 171 AND Y = 21 else
"000000000000" when X = 172 AND Y = 21 else
"000000000000" when X = 173 AND Y = 21 else
"000000000000" when X = 174 AND Y = 21 else
"000000000000" when X = 175 AND Y = 21 else
"000000000000" when X = 176 AND Y = 21 else
"000000000000" when X = 177 AND Y = 21 else
"000000000000" when X = 178 AND Y = 21 else
"000000000000" when X = 179 AND Y = 21 else
"000000000000" when X = 180 AND Y = 21 else
"000000000000" when X = 181 AND Y = 21 else
"000000000000" when X = 182 AND Y = 21 else
"000000000000" when X = 183 AND Y = 21 else
"000000000000" when X = 184 AND Y = 21 else
"000000000000" when X = 185 AND Y = 21 else
"000000000000" when X = 186 AND Y = 21 else
"000000000000" when X = 187 AND Y = 21 else
"000000000000" when X = 188 AND Y = 21 else
"000000000000" when X = 189 AND Y = 21 else
"000000000000" when X = 190 AND Y = 21 else
"000000000000" when X = 191 AND Y = 21 else
"000000000000" when X = 192 AND Y = 21 else
"000000000000" when X = 193 AND Y = 21 else
"000000000000" when X = 194 AND Y = 21 else
"000000000000" when X = 195 AND Y = 21 else
"000000000000" when X = 196 AND Y = 21 else
"000000000000" when X = 197 AND Y = 21 else
"000000000000" when X = 198 AND Y = 21 else
"000000000000" when X = 199 AND Y = 21 else
"000000000000" when X = 200 AND Y = 21 else
"000000000000" when X = 201 AND Y = 21 else
"000000000000" when X = 202 AND Y = 21 else
"000000000000" when X = 203 AND Y = 21 else
"000000000000" when X = 204 AND Y = 21 else
"000000000000" when X = 205 AND Y = 21 else
"000000000000" when X = 206 AND Y = 21 else
"000000000000" when X = 207 AND Y = 21 else
"000000000000" when X = 208 AND Y = 21 else
"000000000000" when X = 209 AND Y = 21 else
"000000000000" when X = 210 AND Y = 21 else
"000000000000" when X = 211 AND Y = 21 else
"000000000000" when X = 212 AND Y = 21 else
"000000000000" when X = 213 AND Y = 21 else
"000000000000" when X = 214 AND Y = 21 else
"000000000000" when X = 215 AND Y = 21 else
"000000000000" when X = 216 AND Y = 21 else
"000000000000" when X = 217 AND Y = 21 else
"000000000000" when X = 218 AND Y = 21 else
"000000000000" when X = 219 AND Y = 21 else
"000000000000" when X = 220 AND Y = 21 else
"000000000000" when X = 221 AND Y = 21 else
"000000000000" when X = 222 AND Y = 21 else
"000000000000" when X = 223 AND Y = 21 else
"000000000000" when X = 224 AND Y = 21 else
"000000000000" when X = 225 AND Y = 21 else
"000000000000" when X = 226 AND Y = 21 else
"000000000000" when X = 227 AND Y = 21 else
"000000000000" when X = 228 AND Y = 21 else
"000000000000" when X = 229 AND Y = 21 else
"000000000000" when X = 230 AND Y = 21 else
"000000000000" when X = 231 AND Y = 21 else
"000000000000" when X = 232 AND Y = 21 else
"000000000000" when X = 233 AND Y = 21 else
"000000000000" when X = 234 AND Y = 21 else
"000000000000" when X = 235 AND Y = 21 else
"000000000000" when X = 236 AND Y = 21 else
"000000000000" when X = 237 AND Y = 21 else
"000000000000" when X = 238 AND Y = 21 else
"000000000000" when X = 239 AND Y = 21 else
"000000000000" when X = 240 AND Y = 21 else
"000000000000" when X = 241 AND Y = 21 else
"000000000000" when X = 242 AND Y = 21 else
"000000000000" when X = 243 AND Y = 21 else
"000000000000" when X = 244 AND Y = 21 else
"000000000000" when X = 245 AND Y = 21 else
"000000000000" when X = 246 AND Y = 21 else
"000000000000" when X = 247 AND Y = 21 else
"000000000000" when X = 248 AND Y = 21 else
"000000000000" when X = 249 AND Y = 21 else
"000000000000" when X = 250 AND Y = 21 else
"000000000000" when X = 251 AND Y = 21 else
"000000000000" when X = 252 AND Y = 21 else
"000000000000" when X = 253 AND Y = 21 else
"000000000000" when X = 254 AND Y = 21 else
"000000000000" when X = 255 AND Y = 21 else
"000000000000" when X = 256 AND Y = 21 else
"000000000000" when X = 257 AND Y = 21 else
"000000000000" when X = 258 AND Y = 21 else
"000000000000" when X = 259 AND Y = 21 else
"000000000000" when X = 260 AND Y = 21 else
"000000000000" when X = 261 AND Y = 21 else
"000000000000" when X = 262 AND Y = 21 else
"000000000000" when X = 263 AND Y = 21 else
"000000000000" when X = 264 AND Y = 21 else
"000000000000" when X = 265 AND Y = 21 else
"000000000000" when X = 266 AND Y = 21 else
"000000000000" when X = 267 AND Y = 21 else
"000000000000" when X = 268 AND Y = 21 else
"000000000000" when X = 269 AND Y = 21 else
"000000000000" when X = 270 AND Y = 21 else
"000000000000" when X = 271 AND Y = 21 else
"000000000000" when X = 272 AND Y = 21 else
"000000000000" when X = 273 AND Y = 21 else
"000000000000" when X = 274 AND Y = 21 else
"000000000000" when X = 275 AND Y = 21 else
"000000000000" when X = 276 AND Y = 21 else
"000000000000" when X = 277 AND Y = 21 else
"000000000000" when X = 278 AND Y = 21 else
"000000000000" when X = 279 AND Y = 21 else
"000000000000" when X = 280 AND Y = 21 else
"000000000000" when X = 281 AND Y = 21 else
"000000000000" when X = 282 AND Y = 21 else
"000000000000" when X = 283 AND Y = 21 else
"000000000000" when X = 284 AND Y = 21 else
"000000000000" when X = 285 AND Y = 21 else
"000000000000" when X = 286 AND Y = 21 else
"000000000000" when X = 287 AND Y = 21 else
"000000000000" when X = 288 AND Y = 21 else
"000000000000" when X = 289 AND Y = 21 else
"000000000000" when X = 290 AND Y = 21 else
"000000000000" when X = 291 AND Y = 21 else
"000000000000" when X = 292 AND Y = 21 else
"000000000000" when X = 293 AND Y = 21 else
"000000000000" when X = 294 AND Y = 21 else
"000000000000" when X = 295 AND Y = 21 else
"000000000000" when X = 296 AND Y = 21 else
"000000000000" when X = 297 AND Y = 21 else
"000000000000" when X = 298 AND Y = 21 else
"000000000000" when X = 299 AND Y = 21 else
"000000000000" when X = 300 AND Y = 21 else
"000000000000" when X = 301 AND Y = 21 else
"000000000000" when X = 302 AND Y = 21 else
"000000000000" when X = 303 AND Y = 21 else
"000000000000" when X = 304 AND Y = 21 else
"000000000000" when X = 305 AND Y = 21 else
"000000000000" when X = 306 AND Y = 21 else
"000000000000" when X = 307 AND Y = 21 else
"000000000000" when X = 308 AND Y = 21 else
"000000000000" when X = 309 AND Y = 21 else
"000000000000" when X = 310 AND Y = 21 else
"000000000000" when X = 311 AND Y = 21 else
"000000000000" when X = 312 AND Y = 21 else
"000000000000" when X = 313 AND Y = 21 else
"000000000000" when X = 314 AND Y = 21 else
"000000000000" when X = 315 AND Y = 21 else
"000000000000" when X = 316 AND Y = 21 else
"000000000000" when X = 317 AND Y = 21 else
"000000000000" when X = 318 AND Y = 21 else
"000000000000" when X = 319 AND Y = 21 else
"000000000000" when X = 320 AND Y = 21 else
"000000000000" when X = 321 AND Y = 21 else
"000000000000" when X = 322 AND Y = 21 else
"000000000000" when X = 323 AND Y = 21 else
"000000000000" when X = 324 AND Y = 21 else
"000000000000" when X = 0 AND Y = 22 else
"000000000000" when X = 1 AND Y = 22 else
"000000000000" when X = 2 AND Y = 22 else
"000000000000" when X = 3 AND Y = 22 else
"000000000000" when X = 4 AND Y = 22 else
"000000000000" when X = 5 AND Y = 22 else
"000000000000" when X = 6 AND Y = 22 else
"000000000000" when X = 7 AND Y = 22 else
"000000000000" when X = 8 AND Y = 22 else
"000000000000" when X = 9 AND Y = 22 else
"000000000000" when X = 10 AND Y = 22 else
"000000000000" when X = 11 AND Y = 22 else
"000000000000" when X = 12 AND Y = 22 else
"000000000000" when X = 13 AND Y = 22 else
"000000000000" when X = 14 AND Y = 22 else
"000000000000" when X = 15 AND Y = 22 else
"000000000000" when X = 16 AND Y = 22 else
"000000000000" when X = 17 AND Y = 22 else
"000000000000" when X = 18 AND Y = 22 else
"000000000000" when X = 19 AND Y = 22 else
"000000000000" when X = 20 AND Y = 22 else
"000000000000" when X = 21 AND Y = 22 else
"000000000000" when X = 22 AND Y = 22 else
"000000000000" when X = 23 AND Y = 22 else
"000000000000" when X = 24 AND Y = 22 else
"000000000000" when X = 25 AND Y = 22 else
"000000000000" when X = 26 AND Y = 22 else
"000000000000" when X = 27 AND Y = 22 else
"000000000000" when X = 28 AND Y = 22 else
"000000000000" when X = 29 AND Y = 22 else
"000000000000" when X = 30 AND Y = 22 else
"000000000000" when X = 31 AND Y = 22 else
"000000000000" when X = 32 AND Y = 22 else
"000000000000" when X = 33 AND Y = 22 else
"000000000000" when X = 34 AND Y = 22 else
"000000000000" when X = 35 AND Y = 22 else
"000000000000" when X = 36 AND Y = 22 else
"000000000000" when X = 37 AND Y = 22 else
"000000000000" when X = 38 AND Y = 22 else
"000000000000" when X = 39 AND Y = 22 else
"100010011101" when X = 40 AND Y = 22 else
"100010011101" when X = 41 AND Y = 22 else
"100010011101" when X = 42 AND Y = 22 else
"100010011101" when X = 43 AND Y = 22 else
"100010011101" when X = 44 AND Y = 22 else
"100010011101" when X = 45 AND Y = 22 else
"100010011101" when X = 46 AND Y = 22 else
"100010011101" when X = 47 AND Y = 22 else
"100010011101" when X = 48 AND Y = 22 else
"100010011101" when X = 49 AND Y = 22 else
"110111011111" when X = 50 AND Y = 22 else
"110111011111" when X = 51 AND Y = 22 else
"110111011111" when X = 52 AND Y = 22 else
"110111011111" when X = 53 AND Y = 22 else
"110111011111" when X = 54 AND Y = 22 else
"110111011111" when X = 55 AND Y = 22 else
"110111011111" when X = 56 AND Y = 22 else
"110111011111" when X = 57 AND Y = 22 else
"110111011111" when X = 58 AND Y = 22 else
"110111011111" when X = 59 AND Y = 22 else
"111111111111" when X = 60 AND Y = 22 else
"111111111111" when X = 61 AND Y = 22 else
"111111111111" when X = 62 AND Y = 22 else
"111111111111" when X = 63 AND Y = 22 else
"111111111111" when X = 64 AND Y = 22 else
"111111111111" when X = 65 AND Y = 22 else
"111111111111" when X = 66 AND Y = 22 else
"111111111111" when X = 67 AND Y = 22 else
"111111111111" when X = 68 AND Y = 22 else
"111111111111" when X = 69 AND Y = 22 else
"111111111111" when X = 70 AND Y = 22 else
"111111111111" when X = 71 AND Y = 22 else
"111111111111" when X = 72 AND Y = 22 else
"111111111111" when X = 73 AND Y = 22 else
"111111111111" when X = 74 AND Y = 22 else
"111111111111" when X = 75 AND Y = 22 else
"111111111111" when X = 76 AND Y = 22 else
"111111111111" when X = 77 AND Y = 22 else
"111111111111" when X = 78 AND Y = 22 else
"111111111111" when X = 79 AND Y = 22 else
"111111111111" when X = 80 AND Y = 22 else
"111111111111" when X = 81 AND Y = 22 else
"111111111111" when X = 82 AND Y = 22 else
"111111111111" when X = 83 AND Y = 22 else
"111111111111" when X = 84 AND Y = 22 else
"111111111111" when X = 85 AND Y = 22 else
"111111111111" when X = 86 AND Y = 22 else
"111111111111" when X = 87 AND Y = 22 else
"111111111111" when X = 88 AND Y = 22 else
"111111111111" when X = 89 AND Y = 22 else
"111111111111" when X = 90 AND Y = 22 else
"111111111111" when X = 91 AND Y = 22 else
"111111111111" when X = 92 AND Y = 22 else
"111111111111" when X = 93 AND Y = 22 else
"111111111111" when X = 94 AND Y = 22 else
"111111111111" when X = 95 AND Y = 22 else
"111111111111" when X = 96 AND Y = 22 else
"111111111111" when X = 97 AND Y = 22 else
"111111111111" when X = 98 AND Y = 22 else
"111111111111" when X = 99 AND Y = 22 else
"111111111111" when X = 100 AND Y = 22 else
"111111111111" when X = 101 AND Y = 22 else
"111111111111" when X = 102 AND Y = 22 else
"111111111111" when X = 103 AND Y = 22 else
"111111111111" when X = 104 AND Y = 22 else
"111111111111" when X = 105 AND Y = 22 else
"111111111111" when X = 106 AND Y = 22 else
"111111111111" when X = 107 AND Y = 22 else
"111111111111" when X = 108 AND Y = 22 else
"111111111111" when X = 109 AND Y = 22 else
"111111111111" when X = 110 AND Y = 22 else
"111111111111" when X = 111 AND Y = 22 else
"111111111111" when X = 112 AND Y = 22 else
"111111111111" when X = 113 AND Y = 22 else
"111111111111" when X = 114 AND Y = 22 else
"111111111111" when X = 115 AND Y = 22 else
"111111111111" when X = 116 AND Y = 22 else
"111111111111" when X = 117 AND Y = 22 else
"111111111111" when X = 118 AND Y = 22 else
"111111111111" when X = 119 AND Y = 22 else
"111111111111" when X = 120 AND Y = 22 else
"111111111111" when X = 121 AND Y = 22 else
"111111111111" when X = 122 AND Y = 22 else
"111111111111" when X = 123 AND Y = 22 else
"111111111111" when X = 124 AND Y = 22 else
"111111111111" when X = 125 AND Y = 22 else
"111111111111" when X = 126 AND Y = 22 else
"111111111111" when X = 127 AND Y = 22 else
"111111111111" when X = 128 AND Y = 22 else
"111111111111" when X = 129 AND Y = 22 else
"111111111111" when X = 130 AND Y = 22 else
"111111111111" when X = 131 AND Y = 22 else
"111111111111" when X = 132 AND Y = 22 else
"111111111111" when X = 133 AND Y = 22 else
"111111111111" when X = 134 AND Y = 22 else
"111111111111" when X = 135 AND Y = 22 else
"111111111111" when X = 136 AND Y = 22 else
"111111111111" when X = 137 AND Y = 22 else
"111111111111" when X = 138 AND Y = 22 else
"111111111111" when X = 139 AND Y = 22 else
"111111111111" when X = 140 AND Y = 22 else
"111111111111" when X = 141 AND Y = 22 else
"111111111111" when X = 142 AND Y = 22 else
"111111111111" when X = 143 AND Y = 22 else
"111111111111" when X = 144 AND Y = 22 else
"111111111111" when X = 145 AND Y = 22 else
"111111111111" when X = 146 AND Y = 22 else
"111111111111" when X = 147 AND Y = 22 else
"111111111111" when X = 148 AND Y = 22 else
"111111111111" when X = 149 AND Y = 22 else
"111111111111" when X = 150 AND Y = 22 else
"111111111111" when X = 151 AND Y = 22 else
"111111111111" when X = 152 AND Y = 22 else
"111111111111" when X = 153 AND Y = 22 else
"111111111111" when X = 154 AND Y = 22 else
"000000000000" when X = 155 AND Y = 22 else
"000000000000" when X = 156 AND Y = 22 else
"000000000000" when X = 157 AND Y = 22 else
"000000000000" when X = 158 AND Y = 22 else
"000000000000" when X = 159 AND Y = 22 else
"000000000000" when X = 160 AND Y = 22 else
"000000000000" when X = 161 AND Y = 22 else
"000000000000" when X = 162 AND Y = 22 else
"000000000000" when X = 163 AND Y = 22 else
"000000000000" when X = 164 AND Y = 22 else
"000000000000" when X = 165 AND Y = 22 else
"000000000000" when X = 166 AND Y = 22 else
"000000000000" when X = 167 AND Y = 22 else
"000000000000" when X = 168 AND Y = 22 else
"000000000000" when X = 169 AND Y = 22 else
"000000000000" when X = 170 AND Y = 22 else
"000000000000" when X = 171 AND Y = 22 else
"000000000000" when X = 172 AND Y = 22 else
"000000000000" when X = 173 AND Y = 22 else
"000000000000" when X = 174 AND Y = 22 else
"000000000000" when X = 175 AND Y = 22 else
"000000000000" when X = 176 AND Y = 22 else
"000000000000" when X = 177 AND Y = 22 else
"000000000000" when X = 178 AND Y = 22 else
"000000000000" when X = 179 AND Y = 22 else
"000000000000" when X = 180 AND Y = 22 else
"000000000000" when X = 181 AND Y = 22 else
"000000000000" when X = 182 AND Y = 22 else
"000000000000" when X = 183 AND Y = 22 else
"000000000000" when X = 184 AND Y = 22 else
"000000000000" when X = 185 AND Y = 22 else
"000000000000" when X = 186 AND Y = 22 else
"000000000000" when X = 187 AND Y = 22 else
"000000000000" when X = 188 AND Y = 22 else
"000000000000" when X = 189 AND Y = 22 else
"000000000000" when X = 190 AND Y = 22 else
"000000000000" when X = 191 AND Y = 22 else
"000000000000" when X = 192 AND Y = 22 else
"000000000000" when X = 193 AND Y = 22 else
"000000000000" when X = 194 AND Y = 22 else
"000000000000" when X = 195 AND Y = 22 else
"000000000000" when X = 196 AND Y = 22 else
"000000000000" when X = 197 AND Y = 22 else
"000000000000" when X = 198 AND Y = 22 else
"000000000000" when X = 199 AND Y = 22 else
"000000000000" when X = 200 AND Y = 22 else
"000000000000" when X = 201 AND Y = 22 else
"000000000000" when X = 202 AND Y = 22 else
"000000000000" when X = 203 AND Y = 22 else
"000000000000" when X = 204 AND Y = 22 else
"000000000000" when X = 205 AND Y = 22 else
"000000000000" when X = 206 AND Y = 22 else
"000000000000" when X = 207 AND Y = 22 else
"000000000000" when X = 208 AND Y = 22 else
"000000000000" when X = 209 AND Y = 22 else
"000000000000" when X = 210 AND Y = 22 else
"000000000000" when X = 211 AND Y = 22 else
"000000000000" when X = 212 AND Y = 22 else
"000000000000" when X = 213 AND Y = 22 else
"000000000000" when X = 214 AND Y = 22 else
"000000000000" when X = 215 AND Y = 22 else
"000000000000" when X = 216 AND Y = 22 else
"000000000000" when X = 217 AND Y = 22 else
"000000000000" when X = 218 AND Y = 22 else
"000000000000" when X = 219 AND Y = 22 else
"000000000000" when X = 220 AND Y = 22 else
"000000000000" when X = 221 AND Y = 22 else
"000000000000" when X = 222 AND Y = 22 else
"000000000000" when X = 223 AND Y = 22 else
"000000000000" when X = 224 AND Y = 22 else
"000000000000" when X = 225 AND Y = 22 else
"000000000000" when X = 226 AND Y = 22 else
"000000000000" when X = 227 AND Y = 22 else
"000000000000" when X = 228 AND Y = 22 else
"000000000000" when X = 229 AND Y = 22 else
"000000000000" when X = 230 AND Y = 22 else
"000000000000" when X = 231 AND Y = 22 else
"000000000000" when X = 232 AND Y = 22 else
"000000000000" when X = 233 AND Y = 22 else
"000000000000" when X = 234 AND Y = 22 else
"000000000000" when X = 235 AND Y = 22 else
"000000000000" when X = 236 AND Y = 22 else
"000000000000" when X = 237 AND Y = 22 else
"000000000000" when X = 238 AND Y = 22 else
"000000000000" when X = 239 AND Y = 22 else
"000000000000" when X = 240 AND Y = 22 else
"000000000000" when X = 241 AND Y = 22 else
"000000000000" when X = 242 AND Y = 22 else
"000000000000" when X = 243 AND Y = 22 else
"000000000000" when X = 244 AND Y = 22 else
"000000000000" when X = 245 AND Y = 22 else
"000000000000" when X = 246 AND Y = 22 else
"000000000000" when X = 247 AND Y = 22 else
"000000000000" when X = 248 AND Y = 22 else
"000000000000" when X = 249 AND Y = 22 else
"000000000000" when X = 250 AND Y = 22 else
"000000000000" when X = 251 AND Y = 22 else
"000000000000" when X = 252 AND Y = 22 else
"000000000000" when X = 253 AND Y = 22 else
"000000000000" when X = 254 AND Y = 22 else
"000000000000" when X = 255 AND Y = 22 else
"000000000000" when X = 256 AND Y = 22 else
"000000000000" when X = 257 AND Y = 22 else
"000000000000" when X = 258 AND Y = 22 else
"000000000000" when X = 259 AND Y = 22 else
"000000000000" when X = 260 AND Y = 22 else
"000000000000" when X = 261 AND Y = 22 else
"000000000000" when X = 262 AND Y = 22 else
"000000000000" when X = 263 AND Y = 22 else
"000000000000" when X = 264 AND Y = 22 else
"000000000000" when X = 265 AND Y = 22 else
"000000000000" when X = 266 AND Y = 22 else
"000000000000" when X = 267 AND Y = 22 else
"000000000000" when X = 268 AND Y = 22 else
"000000000000" when X = 269 AND Y = 22 else
"000000000000" when X = 270 AND Y = 22 else
"000000000000" when X = 271 AND Y = 22 else
"000000000000" when X = 272 AND Y = 22 else
"000000000000" when X = 273 AND Y = 22 else
"000000000000" when X = 274 AND Y = 22 else
"000000000000" when X = 275 AND Y = 22 else
"000000000000" when X = 276 AND Y = 22 else
"000000000000" when X = 277 AND Y = 22 else
"000000000000" when X = 278 AND Y = 22 else
"000000000000" when X = 279 AND Y = 22 else
"000000000000" when X = 280 AND Y = 22 else
"000000000000" when X = 281 AND Y = 22 else
"000000000000" when X = 282 AND Y = 22 else
"000000000000" when X = 283 AND Y = 22 else
"000000000000" when X = 284 AND Y = 22 else
"000000000000" when X = 285 AND Y = 22 else
"000000000000" when X = 286 AND Y = 22 else
"000000000000" when X = 287 AND Y = 22 else
"000000000000" when X = 288 AND Y = 22 else
"000000000000" when X = 289 AND Y = 22 else
"000000000000" when X = 290 AND Y = 22 else
"000000000000" when X = 291 AND Y = 22 else
"000000000000" when X = 292 AND Y = 22 else
"000000000000" when X = 293 AND Y = 22 else
"000000000000" when X = 294 AND Y = 22 else
"000000000000" when X = 295 AND Y = 22 else
"000000000000" when X = 296 AND Y = 22 else
"000000000000" when X = 297 AND Y = 22 else
"000000000000" when X = 298 AND Y = 22 else
"000000000000" when X = 299 AND Y = 22 else
"000000000000" when X = 300 AND Y = 22 else
"000000000000" when X = 301 AND Y = 22 else
"000000000000" when X = 302 AND Y = 22 else
"000000000000" when X = 303 AND Y = 22 else
"000000000000" when X = 304 AND Y = 22 else
"000000000000" when X = 305 AND Y = 22 else
"000000000000" when X = 306 AND Y = 22 else
"000000000000" when X = 307 AND Y = 22 else
"000000000000" when X = 308 AND Y = 22 else
"000000000000" when X = 309 AND Y = 22 else
"000000000000" when X = 310 AND Y = 22 else
"000000000000" when X = 311 AND Y = 22 else
"000000000000" when X = 312 AND Y = 22 else
"000000000000" when X = 313 AND Y = 22 else
"000000000000" when X = 314 AND Y = 22 else
"000000000000" when X = 315 AND Y = 22 else
"000000000000" when X = 316 AND Y = 22 else
"000000000000" when X = 317 AND Y = 22 else
"000000000000" when X = 318 AND Y = 22 else
"000000000000" when X = 319 AND Y = 22 else
"000000000000" when X = 320 AND Y = 22 else
"000000000000" when X = 321 AND Y = 22 else
"000000000000" when X = 322 AND Y = 22 else
"000000000000" when X = 323 AND Y = 22 else
"000000000000" when X = 324 AND Y = 22 else
"000000000000" when X = 0 AND Y = 23 else
"000000000000" when X = 1 AND Y = 23 else
"000000000000" when X = 2 AND Y = 23 else
"000000000000" when X = 3 AND Y = 23 else
"000000000000" when X = 4 AND Y = 23 else
"000000000000" when X = 5 AND Y = 23 else
"000000000000" when X = 6 AND Y = 23 else
"000000000000" when X = 7 AND Y = 23 else
"000000000000" when X = 8 AND Y = 23 else
"000000000000" when X = 9 AND Y = 23 else
"000000000000" when X = 10 AND Y = 23 else
"000000000000" when X = 11 AND Y = 23 else
"000000000000" when X = 12 AND Y = 23 else
"000000000000" when X = 13 AND Y = 23 else
"000000000000" when X = 14 AND Y = 23 else
"000000000000" when X = 15 AND Y = 23 else
"000000000000" when X = 16 AND Y = 23 else
"000000000000" when X = 17 AND Y = 23 else
"000000000000" when X = 18 AND Y = 23 else
"000000000000" when X = 19 AND Y = 23 else
"000000000000" when X = 20 AND Y = 23 else
"000000000000" when X = 21 AND Y = 23 else
"000000000000" when X = 22 AND Y = 23 else
"000000000000" when X = 23 AND Y = 23 else
"000000000000" when X = 24 AND Y = 23 else
"000000000000" when X = 25 AND Y = 23 else
"000000000000" when X = 26 AND Y = 23 else
"000000000000" when X = 27 AND Y = 23 else
"000000000000" when X = 28 AND Y = 23 else
"000000000000" when X = 29 AND Y = 23 else
"000000000000" when X = 30 AND Y = 23 else
"000000000000" when X = 31 AND Y = 23 else
"000000000000" when X = 32 AND Y = 23 else
"000000000000" when X = 33 AND Y = 23 else
"000000000000" when X = 34 AND Y = 23 else
"000000000000" when X = 35 AND Y = 23 else
"000000000000" when X = 36 AND Y = 23 else
"000000000000" when X = 37 AND Y = 23 else
"000000000000" when X = 38 AND Y = 23 else
"000000000000" when X = 39 AND Y = 23 else
"100010011101" when X = 40 AND Y = 23 else
"100010011101" when X = 41 AND Y = 23 else
"100010011101" when X = 42 AND Y = 23 else
"100010011101" when X = 43 AND Y = 23 else
"100010011101" when X = 44 AND Y = 23 else
"100010011101" when X = 45 AND Y = 23 else
"100010011101" when X = 46 AND Y = 23 else
"100010011101" when X = 47 AND Y = 23 else
"100010011101" when X = 48 AND Y = 23 else
"100010011101" when X = 49 AND Y = 23 else
"110111011111" when X = 50 AND Y = 23 else
"110111011111" when X = 51 AND Y = 23 else
"110111011111" when X = 52 AND Y = 23 else
"110111011111" when X = 53 AND Y = 23 else
"110111011111" when X = 54 AND Y = 23 else
"110111011111" when X = 55 AND Y = 23 else
"110111011111" when X = 56 AND Y = 23 else
"110111011111" when X = 57 AND Y = 23 else
"110111011111" when X = 58 AND Y = 23 else
"110111011111" when X = 59 AND Y = 23 else
"111111111111" when X = 60 AND Y = 23 else
"111111111111" when X = 61 AND Y = 23 else
"111111111111" when X = 62 AND Y = 23 else
"111111111111" when X = 63 AND Y = 23 else
"111111111111" when X = 64 AND Y = 23 else
"111111111111" when X = 65 AND Y = 23 else
"111111111111" when X = 66 AND Y = 23 else
"111111111111" when X = 67 AND Y = 23 else
"111111111111" when X = 68 AND Y = 23 else
"111111111111" when X = 69 AND Y = 23 else
"111111111111" when X = 70 AND Y = 23 else
"111111111111" when X = 71 AND Y = 23 else
"111111111111" when X = 72 AND Y = 23 else
"111111111111" when X = 73 AND Y = 23 else
"111111111111" when X = 74 AND Y = 23 else
"111111111111" when X = 75 AND Y = 23 else
"111111111111" when X = 76 AND Y = 23 else
"111111111111" when X = 77 AND Y = 23 else
"111111111111" when X = 78 AND Y = 23 else
"111111111111" when X = 79 AND Y = 23 else
"111111111111" when X = 80 AND Y = 23 else
"111111111111" when X = 81 AND Y = 23 else
"111111111111" when X = 82 AND Y = 23 else
"111111111111" when X = 83 AND Y = 23 else
"111111111111" when X = 84 AND Y = 23 else
"111111111111" when X = 85 AND Y = 23 else
"111111111111" when X = 86 AND Y = 23 else
"111111111111" when X = 87 AND Y = 23 else
"111111111111" when X = 88 AND Y = 23 else
"111111111111" when X = 89 AND Y = 23 else
"111111111111" when X = 90 AND Y = 23 else
"111111111111" when X = 91 AND Y = 23 else
"111111111111" when X = 92 AND Y = 23 else
"111111111111" when X = 93 AND Y = 23 else
"111111111111" when X = 94 AND Y = 23 else
"111111111111" when X = 95 AND Y = 23 else
"111111111111" when X = 96 AND Y = 23 else
"111111111111" when X = 97 AND Y = 23 else
"111111111111" when X = 98 AND Y = 23 else
"111111111111" when X = 99 AND Y = 23 else
"111111111111" when X = 100 AND Y = 23 else
"111111111111" when X = 101 AND Y = 23 else
"111111111111" when X = 102 AND Y = 23 else
"111111111111" when X = 103 AND Y = 23 else
"111111111111" when X = 104 AND Y = 23 else
"111111111111" when X = 105 AND Y = 23 else
"111111111111" when X = 106 AND Y = 23 else
"111111111111" when X = 107 AND Y = 23 else
"111111111111" when X = 108 AND Y = 23 else
"111111111111" when X = 109 AND Y = 23 else
"111111111111" when X = 110 AND Y = 23 else
"111111111111" when X = 111 AND Y = 23 else
"111111111111" when X = 112 AND Y = 23 else
"111111111111" when X = 113 AND Y = 23 else
"111111111111" when X = 114 AND Y = 23 else
"111111111111" when X = 115 AND Y = 23 else
"111111111111" when X = 116 AND Y = 23 else
"111111111111" when X = 117 AND Y = 23 else
"111111111111" when X = 118 AND Y = 23 else
"111111111111" when X = 119 AND Y = 23 else
"111111111111" when X = 120 AND Y = 23 else
"111111111111" when X = 121 AND Y = 23 else
"111111111111" when X = 122 AND Y = 23 else
"111111111111" when X = 123 AND Y = 23 else
"111111111111" when X = 124 AND Y = 23 else
"111111111111" when X = 125 AND Y = 23 else
"111111111111" when X = 126 AND Y = 23 else
"111111111111" when X = 127 AND Y = 23 else
"111111111111" when X = 128 AND Y = 23 else
"111111111111" when X = 129 AND Y = 23 else
"111111111111" when X = 130 AND Y = 23 else
"111111111111" when X = 131 AND Y = 23 else
"111111111111" when X = 132 AND Y = 23 else
"111111111111" when X = 133 AND Y = 23 else
"111111111111" when X = 134 AND Y = 23 else
"111111111111" when X = 135 AND Y = 23 else
"111111111111" when X = 136 AND Y = 23 else
"111111111111" when X = 137 AND Y = 23 else
"111111111111" when X = 138 AND Y = 23 else
"111111111111" when X = 139 AND Y = 23 else
"111111111111" when X = 140 AND Y = 23 else
"111111111111" when X = 141 AND Y = 23 else
"111111111111" when X = 142 AND Y = 23 else
"111111111111" when X = 143 AND Y = 23 else
"111111111111" when X = 144 AND Y = 23 else
"111111111111" when X = 145 AND Y = 23 else
"111111111111" when X = 146 AND Y = 23 else
"111111111111" when X = 147 AND Y = 23 else
"111111111111" when X = 148 AND Y = 23 else
"111111111111" when X = 149 AND Y = 23 else
"111111111111" when X = 150 AND Y = 23 else
"111111111111" when X = 151 AND Y = 23 else
"111111111111" when X = 152 AND Y = 23 else
"111111111111" when X = 153 AND Y = 23 else
"111111111111" when X = 154 AND Y = 23 else
"000000000000" when X = 155 AND Y = 23 else
"000000000000" when X = 156 AND Y = 23 else
"000000000000" when X = 157 AND Y = 23 else
"000000000000" when X = 158 AND Y = 23 else
"000000000000" when X = 159 AND Y = 23 else
"000000000000" when X = 160 AND Y = 23 else
"000000000000" when X = 161 AND Y = 23 else
"000000000000" when X = 162 AND Y = 23 else
"000000000000" when X = 163 AND Y = 23 else
"000000000000" when X = 164 AND Y = 23 else
"000000000000" when X = 165 AND Y = 23 else
"000000000000" when X = 166 AND Y = 23 else
"000000000000" when X = 167 AND Y = 23 else
"000000000000" when X = 168 AND Y = 23 else
"000000000000" when X = 169 AND Y = 23 else
"000000000000" when X = 170 AND Y = 23 else
"000000000000" when X = 171 AND Y = 23 else
"000000000000" when X = 172 AND Y = 23 else
"000000000000" when X = 173 AND Y = 23 else
"000000000000" when X = 174 AND Y = 23 else
"000000000000" when X = 175 AND Y = 23 else
"000000000000" when X = 176 AND Y = 23 else
"000000000000" when X = 177 AND Y = 23 else
"000000000000" when X = 178 AND Y = 23 else
"000000000000" when X = 179 AND Y = 23 else
"000000000000" when X = 180 AND Y = 23 else
"000000000000" when X = 181 AND Y = 23 else
"000000000000" when X = 182 AND Y = 23 else
"000000000000" when X = 183 AND Y = 23 else
"000000000000" when X = 184 AND Y = 23 else
"000000000000" when X = 185 AND Y = 23 else
"000000000000" when X = 186 AND Y = 23 else
"000000000000" when X = 187 AND Y = 23 else
"000000000000" when X = 188 AND Y = 23 else
"000000000000" when X = 189 AND Y = 23 else
"000000000000" when X = 190 AND Y = 23 else
"000000000000" when X = 191 AND Y = 23 else
"000000000000" when X = 192 AND Y = 23 else
"000000000000" when X = 193 AND Y = 23 else
"000000000000" when X = 194 AND Y = 23 else
"000000000000" when X = 195 AND Y = 23 else
"000000000000" when X = 196 AND Y = 23 else
"000000000000" when X = 197 AND Y = 23 else
"000000000000" when X = 198 AND Y = 23 else
"000000000000" when X = 199 AND Y = 23 else
"000000000000" when X = 200 AND Y = 23 else
"000000000000" when X = 201 AND Y = 23 else
"000000000000" when X = 202 AND Y = 23 else
"000000000000" when X = 203 AND Y = 23 else
"000000000000" when X = 204 AND Y = 23 else
"000000000000" when X = 205 AND Y = 23 else
"000000000000" when X = 206 AND Y = 23 else
"000000000000" when X = 207 AND Y = 23 else
"000000000000" when X = 208 AND Y = 23 else
"000000000000" when X = 209 AND Y = 23 else
"000000000000" when X = 210 AND Y = 23 else
"000000000000" when X = 211 AND Y = 23 else
"000000000000" when X = 212 AND Y = 23 else
"000000000000" when X = 213 AND Y = 23 else
"000000000000" when X = 214 AND Y = 23 else
"000000000000" when X = 215 AND Y = 23 else
"000000000000" when X = 216 AND Y = 23 else
"000000000000" when X = 217 AND Y = 23 else
"000000000000" when X = 218 AND Y = 23 else
"000000000000" when X = 219 AND Y = 23 else
"000000000000" when X = 220 AND Y = 23 else
"000000000000" when X = 221 AND Y = 23 else
"000000000000" when X = 222 AND Y = 23 else
"000000000000" when X = 223 AND Y = 23 else
"000000000000" when X = 224 AND Y = 23 else
"000000000000" when X = 225 AND Y = 23 else
"000000000000" when X = 226 AND Y = 23 else
"000000000000" when X = 227 AND Y = 23 else
"000000000000" when X = 228 AND Y = 23 else
"000000000000" when X = 229 AND Y = 23 else
"000000000000" when X = 230 AND Y = 23 else
"000000000000" when X = 231 AND Y = 23 else
"000000000000" when X = 232 AND Y = 23 else
"000000000000" when X = 233 AND Y = 23 else
"000000000000" when X = 234 AND Y = 23 else
"000000000000" when X = 235 AND Y = 23 else
"000000000000" when X = 236 AND Y = 23 else
"000000000000" when X = 237 AND Y = 23 else
"000000000000" when X = 238 AND Y = 23 else
"000000000000" when X = 239 AND Y = 23 else
"000000000000" when X = 240 AND Y = 23 else
"000000000000" when X = 241 AND Y = 23 else
"000000000000" when X = 242 AND Y = 23 else
"000000000000" when X = 243 AND Y = 23 else
"000000000000" when X = 244 AND Y = 23 else
"000000000000" when X = 245 AND Y = 23 else
"000000000000" when X = 246 AND Y = 23 else
"000000000000" when X = 247 AND Y = 23 else
"000000000000" when X = 248 AND Y = 23 else
"000000000000" when X = 249 AND Y = 23 else
"000000000000" when X = 250 AND Y = 23 else
"000000000000" when X = 251 AND Y = 23 else
"000000000000" when X = 252 AND Y = 23 else
"000000000000" when X = 253 AND Y = 23 else
"000000000000" when X = 254 AND Y = 23 else
"000000000000" when X = 255 AND Y = 23 else
"000000000000" when X = 256 AND Y = 23 else
"000000000000" when X = 257 AND Y = 23 else
"000000000000" when X = 258 AND Y = 23 else
"000000000000" when X = 259 AND Y = 23 else
"000000000000" when X = 260 AND Y = 23 else
"000000000000" when X = 261 AND Y = 23 else
"000000000000" when X = 262 AND Y = 23 else
"000000000000" when X = 263 AND Y = 23 else
"000000000000" when X = 264 AND Y = 23 else
"000000000000" when X = 265 AND Y = 23 else
"000000000000" when X = 266 AND Y = 23 else
"000000000000" when X = 267 AND Y = 23 else
"000000000000" when X = 268 AND Y = 23 else
"000000000000" when X = 269 AND Y = 23 else
"000000000000" when X = 270 AND Y = 23 else
"000000000000" when X = 271 AND Y = 23 else
"000000000000" when X = 272 AND Y = 23 else
"000000000000" when X = 273 AND Y = 23 else
"000000000000" when X = 274 AND Y = 23 else
"000000000000" when X = 275 AND Y = 23 else
"000000000000" when X = 276 AND Y = 23 else
"000000000000" when X = 277 AND Y = 23 else
"000000000000" when X = 278 AND Y = 23 else
"000000000000" when X = 279 AND Y = 23 else
"000000000000" when X = 280 AND Y = 23 else
"000000000000" when X = 281 AND Y = 23 else
"000000000000" when X = 282 AND Y = 23 else
"000000000000" when X = 283 AND Y = 23 else
"000000000000" when X = 284 AND Y = 23 else
"000000000000" when X = 285 AND Y = 23 else
"000000000000" when X = 286 AND Y = 23 else
"000000000000" when X = 287 AND Y = 23 else
"000000000000" when X = 288 AND Y = 23 else
"000000000000" when X = 289 AND Y = 23 else
"000000000000" when X = 290 AND Y = 23 else
"000000000000" when X = 291 AND Y = 23 else
"000000000000" when X = 292 AND Y = 23 else
"000000000000" when X = 293 AND Y = 23 else
"000000000000" when X = 294 AND Y = 23 else
"000000000000" when X = 295 AND Y = 23 else
"000000000000" when X = 296 AND Y = 23 else
"000000000000" when X = 297 AND Y = 23 else
"000000000000" when X = 298 AND Y = 23 else
"000000000000" when X = 299 AND Y = 23 else
"000000000000" when X = 300 AND Y = 23 else
"000000000000" when X = 301 AND Y = 23 else
"000000000000" when X = 302 AND Y = 23 else
"000000000000" when X = 303 AND Y = 23 else
"000000000000" when X = 304 AND Y = 23 else
"000000000000" when X = 305 AND Y = 23 else
"000000000000" when X = 306 AND Y = 23 else
"000000000000" when X = 307 AND Y = 23 else
"000000000000" when X = 308 AND Y = 23 else
"000000000000" when X = 309 AND Y = 23 else
"000000000000" when X = 310 AND Y = 23 else
"000000000000" when X = 311 AND Y = 23 else
"000000000000" when X = 312 AND Y = 23 else
"000000000000" when X = 313 AND Y = 23 else
"000000000000" when X = 314 AND Y = 23 else
"000000000000" when X = 315 AND Y = 23 else
"000000000000" when X = 316 AND Y = 23 else
"000000000000" when X = 317 AND Y = 23 else
"000000000000" when X = 318 AND Y = 23 else
"000000000000" when X = 319 AND Y = 23 else
"000000000000" when X = 320 AND Y = 23 else
"000000000000" when X = 321 AND Y = 23 else
"000000000000" when X = 322 AND Y = 23 else
"000000000000" when X = 323 AND Y = 23 else
"000000000000" when X = 324 AND Y = 23 else
"000000000000" when X = 0 AND Y = 24 else
"000000000000" when X = 1 AND Y = 24 else
"000000000000" when X = 2 AND Y = 24 else
"000000000000" when X = 3 AND Y = 24 else
"000000000000" when X = 4 AND Y = 24 else
"000000000000" when X = 5 AND Y = 24 else
"000000000000" when X = 6 AND Y = 24 else
"000000000000" when X = 7 AND Y = 24 else
"000000000000" when X = 8 AND Y = 24 else
"000000000000" when X = 9 AND Y = 24 else
"000000000000" when X = 10 AND Y = 24 else
"000000000000" when X = 11 AND Y = 24 else
"000000000000" when X = 12 AND Y = 24 else
"000000000000" when X = 13 AND Y = 24 else
"000000000000" when X = 14 AND Y = 24 else
"000000000000" when X = 15 AND Y = 24 else
"000000000000" when X = 16 AND Y = 24 else
"000000000000" when X = 17 AND Y = 24 else
"000000000000" when X = 18 AND Y = 24 else
"000000000000" when X = 19 AND Y = 24 else
"000000000000" when X = 20 AND Y = 24 else
"000000000000" when X = 21 AND Y = 24 else
"000000000000" when X = 22 AND Y = 24 else
"000000000000" when X = 23 AND Y = 24 else
"000000000000" when X = 24 AND Y = 24 else
"000000000000" when X = 25 AND Y = 24 else
"000000000000" when X = 26 AND Y = 24 else
"000000000000" when X = 27 AND Y = 24 else
"000000000000" when X = 28 AND Y = 24 else
"000000000000" when X = 29 AND Y = 24 else
"000000000000" when X = 30 AND Y = 24 else
"000000000000" when X = 31 AND Y = 24 else
"000000000000" when X = 32 AND Y = 24 else
"000000000000" when X = 33 AND Y = 24 else
"000000000000" when X = 34 AND Y = 24 else
"000000000000" when X = 35 AND Y = 24 else
"000000000000" when X = 36 AND Y = 24 else
"000000000000" when X = 37 AND Y = 24 else
"000000000000" when X = 38 AND Y = 24 else
"000000000000" when X = 39 AND Y = 24 else
"100010011101" when X = 40 AND Y = 24 else
"100010011101" when X = 41 AND Y = 24 else
"100010011101" when X = 42 AND Y = 24 else
"100010011101" when X = 43 AND Y = 24 else
"100010011101" when X = 44 AND Y = 24 else
"100010011101" when X = 45 AND Y = 24 else
"100010011101" when X = 46 AND Y = 24 else
"100010011101" when X = 47 AND Y = 24 else
"100010011101" when X = 48 AND Y = 24 else
"100010011101" when X = 49 AND Y = 24 else
"110111011111" when X = 50 AND Y = 24 else
"110111011111" when X = 51 AND Y = 24 else
"110111011111" when X = 52 AND Y = 24 else
"110111011111" when X = 53 AND Y = 24 else
"110111011111" when X = 54 AND Y = 24 else
"110111011111" when X = 55 AND Y = 24 else
"110111011111" when X = 56 AND Y = 24 else
"110111011111" when X = 57 AND Y = 24 else
"110111011111" when X = 58 AND Y = 24 else
"110111011111" when X = 59 AND Y = 24 else
"111111111111" when X = 60 AND Y = 24 else
"111111111111" when X = 61 AND Y = 24 else
"111111111111" when X = 62 AND Y = 24 else
"111111111111" when X = 63 AND Y = 24 else
"111111111111" when X = 64 AND Y = 24 else
"111111111111" when X = 65 AND Y = 24 else
"111111111111" when X = 66 AND Y = 24 else
"111111111111" when X = 67 AND Y = 24 else
"111111111111" when X = 68 AND Y = 24 else
"111111111111" when X = 69 AND Y = 24 else
"111111111111" when X = 70 AND Y = 24 else
"111111111111" when X = 71 AND Y = 24 else
"111111111111" when X = 72 AND Y = 24 else
"111111111111" when X = 73 AND Y = 24 else
"111111111111" when X = 74 AND Y = 24 else
"111111111111" when X = 75 AND Y = 24 else
"111111111111" when X = 76 AND Y = 24 else
"111111111111" when X = 77 AND Y = 24 else
"111111111111" when X = 78 AND Y = 24 else
"111111111111" when X = 79 AND Y = 24 else
"111111111111" when X = 80 AND Y = 24 else
"111111111111" when X = 81 AND Y = 24 else
"111111111111" when X = 82 AND Y = 24 else
"111111111111" when X = 83 AND Y = 24 else
"111111111111" when X = 84 AND Y = 24 else
"111111111111" when X = 85 AND Y = 24 else
"111111111111" when X = 86 AND Y = 24 else
"111111111111" when X = 87 AND Y = 24 else
"111111111111" when X = 88 AND Y = 24 else
"111111111111" when X = 89 AND Y = 24 else
"111111111111" when X = 90 AND Y = 24 else
"111111111111" when X = 91 AND Y = 24 else
"111111111111" when X = 92 AND Y = 24 else
"111111111111" when X = 93 AND Y = 24 else
"111111111111" when X = 94 AND Y = 24 else
"111111111111" when X = 95 AND Y = 24 else
"111111111111" when X = 96 AND Y = 24 else
"111111111111" when X = 97 AND Y = 24 else
"111111111111" when X = 98 AND Y = 24 else
"111111111111" when X = 99 AND Y = 24 else
"111111111111" when X = 100 AND Y = 24 else
"111111111111" when X = 101 AND Y = 24 else
"111111111111" when X = 102 AND Y = 24 else
"111111111111" when X = 103 AND Y = 24 else
"111111111111" when X = 104 AND Y = 24 else
"111111111111" when X = 105 AND Y = 24 else
"111111111111" when X = 106 AND Y = 24 else
"111111111111" when X = 107 AND Y = 24 else
"111111111111" when X = 108 AND Y = 24 else
"111111111111" when X = 109 AND Y = 24 else
"111111111111" when X = 110 AND Y = 24 else
"111111111111" when X = 111 AND Y = 24 else
"111111111111" when X = 112 AND Y = 24 else
"111111111111" when X = 113 AND Y = 24 else
"111111111111" when X = 114 AND Y = 24 else
"111111111111" when X = 115 AND Y = 24 else
"111111111111" when X = 116 AND Y = 24 else
"111111111111" when X = 117 AND Y = 24 else
"111111111111" when X = 118 AND Y = 24 else
"111111111111" when X = 119 AND Y = 24 else
"111111111111" when X = 120 AND Y = 24 else
"111111111111" when X = 121 AND Y = 24 else
"111111111111" when X = 122 AND Y = 24 else
"111111111111" when X = 123 AND Y = 24 else
"111111111111" when X = 124 AND Y = 24 else
"111111111111" when X = 125 AND Y = 24 else
"111111111111" when X = 126 AND Y = 24 else
"111111111111" when X = 127 AND Y = 24 else
"111111111111" when X = 128 AND Y = 24 else
"111111111111" when X = 129 AND Y = 24 else
"111111111111" when X = 130 AND Y = 24 else
"111111111111" when X = 131 AND Y = 24 else
"111111111111" when X = 132 AND Y = 24 else
"111111111111" when X = 133 AND Y = 24 else
"111111111111" when X = 134 AND Y = 24 else
"111111111111" when X = 135 AND Y = 24 else
"111111111111" when X = 136 AND Y = 24 else
"111111111111" when X = 137 AND Y = 24 else
"111111111111" when X = 138 AND Y = 24 else
"111111111111" when X = 139 AND Y = 24 else
"111111111111" when X = 140 AND Y = 24 else
"111111111111" when X = 141 AND Y = 24 else
"111111111111" when X = 142 AND Y = 24 else
"111111111111" when X = 143 AND Y = 24 else
"111111111111" when X = 144 AND Y = 24 else
"111111111111" when X = 145 AND Y = 24 else
"111111111111" when X = 146 AND Y = 24 else
"111111111111" when X = 147 AND Y = 24 else
"111111111111" when X = 148 AND Y = 24 else
"111111111111" when X = 149 AND Y = 24 else
"111111111111" when X = 150 AND Y = 24 else
"111111111111" when X = 151 AND Y = 24 else
"111111111111" when X = 152 AND Y = 24 else
"111111111111" when X = 153 AND Y = 24 else
"111111111111" when X = 154 AND Y = 24 else
"000000000000" when X = 155 AND Y = 24 else
"000000000000" when X = 156 AND Y = 24 else
"000000000000" when X = 157 AND Y = 24 else
"000000000000" when X = 158 AND Y = 24 else
"000000000000" when X = 159 AND Y = 24 else
"000000000000" when X = 160 AND Y = 24 else
"000000000000" when X = 161 AND Y = 24 else
"000000000000" when X = 162 AND Y = 24 else
"000000000000" when X = 163 AND Y = 24 else
"000000000000" when X = 164 AND Y = 24 else
"000000000000" when X = 165 AND Y = 24 else
"000000000000" when X = 166 AND Y = 24 else
"000000000000" when X = 167 AND Y = 24 else
"000000000000" when X = 168 AND Y = 24 else
"000000000000" when X = 169 AND Y = 24 else
"000000000000" when X = 170 AND Y = 24 else
"000000000000" when X = 171 AND Y = 24 else
"000000000000" when X = 172 AND Y = 24 else
"000000000000" when X = 173 AND Y = 24 else
"000000000000" when X = 174 AND Y = 24 else
"000000000000" when X = 175 AND Y = 24 else
"000000000000" when X = 176 AND Y = 24 else
"000000000000" when X = 177 AND Y = 24 else
"000000000000" when X = 178 AND Y = 24 else
"000000000000" when X = 179 AND Y = 24 else
"000000000000" when X = 180 AND Y = 24 else
"000000000000" when X = 181 AND Y = 24 else
"000000000000" when X = 182 AND Y = 24 else
"000000000000" when X = 183 AND Y = 24 else
"000000000000" when X = 184 AND Y = 24 else
"000000000000" when X = 185 AND Y = 24 else
"000000000000" when X = 186 AND Y = 24 else
"000000000000" when X = 187 AND Y = 24 else
"000000000000" when X = 188 AND Y = 24 else
"000000000000" when X = 189 AND Y = 24 else
"000000000000" when X = 190 AND Y = 24 else
"000000000000" when X = 191 AND Y = 24 else
"000000000000" when X = 192 AND Y = 24 else
"000000000000" when X = 193 AND Y = 24 else
"000000000000" when X = 194 AND Y = 24 else
"000000000000" when X = 195 AND Y = 24 else
"000000000000" when X = 196 AND Y = 24 else
"000000000000" when X = 197 AND Y = 24 else
"000000000000" when X = 198 AND Y = 24 else
"000000000000" when X = 199 AND Y = 24 else
"000000000000" when X = 200 AND Y = 24 else
"000000000000" when X = 201 AND Y = 24 else
"000000000000" when X = 202 AND Y = 24 else
"000000000000" when X = 203 AND Y = 24 else
"000000000000" when X = 204 AND Y = 24 else
"000000000000" when X = 205 AND Y = 24 else
"000000000000" when X = 206 AND Y = 24 else
"000000000000" when X = 207 AND Y = 24 else
"000000000000" when X = 208 AND Y = 24 else
"000000000000" when X = 209 AND Y = 24 else
"000000000000" when X = 210 AND Y = 24 else
"000000000000" when X = 211 AND Y = 24 else
"000000000000" when X = 212 AND Y = 24 else
"000000000000" when X = 213 AND Y = 24 else
"000000000000" when X = 214 AND Y = 24 else
"000000000000" when X = 215 AND Y = 24 else
"000000000000" when X = 216 AND Y = 24 else
"000000000000" when X = 217 AND Y = 24 else
"000000000000" when X = 218 AND Y = 24 else
"000000000000" when X = 219 AND Y = 24 else
"000000000000" when X = 220 AND Y = 24 else
"000000000000" when X = 221 AND Y = 24 else
"000000000000" when X = 222 AND Y = 24 else
"000000000000" when X = 223 AND Y = 24 else
"000000000000" when X = 224 AND Y = 24 else
"000000000000" when X = 225 AND Y = 24 else
"000000000000" when X = 226 AND Y = 24 else
"000000000000" when X = 227 AND Y = 24 else
"000000000000" when X = 228 AND Y = 24 else
"000000000000" when X = 229 AND Y = 24 else
"000000000000" when X = 230 AND Y = 24 else
"000000000000" when X = 231 AND Y = 24 else
"000000000000" when X = 232 AND Y = 24 else
"000000000000" when X = 233 AND Y = 24 else
"000000000000" when X = 234 AND Y = 24 else
"000000000000" when X = 235 AND Y = 24 else
"000000000000" when X = 236 AND Y = 24 else
"000000000000" when X = 237 AND Y = 24 else
"000000000000" when X = 238 AND Y = 24 else
"000000000000" when X = 239 AND Y = 24 else
"000000000000" when X = 240 AND Y = 24 else
"000000000000" when X = 241 AND Y = 24 else
"000000000000" when X = 242 AND Y = 24 else
"000000000000" when X = 243 AND Y = 24 else
"000000000000" when X = 244 AND Y = 24 else
"000000000000" when X = 245 AND Y = 24 else
"000000000000" when X = 246 AND Y = 24 else
"000000000000" when X = 247 AND Y = 24 else
"000000000000" when X = 248 AND Y = 24 else
"000000000000" when X = 249 AND Y = 24 else
"000000000000" when X = 250 AND Y = 24 else
"000000000000" when X = 251 AND Y = 24 else
"000000000000" when X = 252 AND Y = 24 else
"000000000000" when X = 253 AND Y = 24 else
"000000000000" when X = 254 AND Y = 24 else
"000000000000" when X = 255 AND Y = 24 else
"000000000000" when X = 256 AND Y = 24 else
"000000000000" when X = 257 AND Y = 24 else
"000000000000" when X = 258 AND Y = 24 else
"000000000000" when X = 259 AND Y = 24 else
"000000000000" when X = 260 AND Y = 24 else
"000000000000" when X = 261 AND Y = 24 else
"000000000000" when X = 262 AND Y = 24 else
"000000000000" when X = 263 AND Y = 24 else
"000000000000" when X = 264 AND Y = 24 else
"000000000000" when X = 265 AND Y = 24 else
"000000000000" when X = 266 AND Y = 24 else
"000000000000" when X = 267 AND Y = 24 else
"000000000000" when X = 268 AND Y = 24 else
"000000000000" when X = 269 AND Y = 24 else
"000000000000" when X = 270 AND Y = 24 else
"000000000000" when X = 271 AND Y = 24 else
"000000000000" when X = 272 AND Y = 24 else
"000000000000" when X = 273 AND Y = 24 else
"000000000000" when X = 274 AND Y = 24 else
"000000000000" when X = 275 AND Y = 24 else
"000000000000" when X = 276 AND Y = 24 else
"000000000000" when X = 277 AND Y = 24 else
"000000000000" when X = 278 AND Y = 24 else
"000000000000" when X = 279 AND Y = 24 else
"000000000000" when X = 280 AND Y = 24 else
"000000000000" when X = 281 AND Y = 24 else
"000000000000" when X = 282 AND Y = 24 else
"000000000000" when X = 283 AND Y = 24 else
"000000000000" when X = 284 AND Y = 24 else
"000000000000" when X = 285 AND Y = 24 else
"000000000000" when X = 286 AND Y = 24 else
"000000000000" when X = 287 AND Y = 24 else
"000000000000" when X = 288 AND Y = 24 else
"000000000000" when X = 289 AND Y = 24 else
"000000000000" when X = 290 AND Y = 24 else
"000000000000" when X = 291 AND Y = 24 else
"000000000000" when X = 292 AND Y = 24 else
"000000000000" when X = 293 AND Y = 24 else
"000000000000" when X = 294 AND Y = 24 else
"000000000000" when X = 295 AND Y = 24 else
"000000000000" when X = 296 AND Y = 24 else
"000000000000" when X = 297 AND Y = 24 else
"000000000000" when X = 298 AND Y = 24 else
"000000000000" when X = 299 AND Y = 24 else
"000000000000" when X = 300 AND Y = 24 else
"000000000000" when X = 301 AND Y = 24 else
"000000000000" when X = 302 AND Y = 24 else
"000000000000" when X = 303 AND Y = 24 else
"000000000000" when X = 304 AND Y = 24 else
"000000000000" when X = 305 AND Y = 24 else
"000000000000" when X = 306 AND Y = 24 else
"000000000000" when X = 307 AND Y = 24 else
"000000000000" when X = 308 AND Y = 24 else
"000000000000" when X = 309 AND Y = 24 else
"000000000000" when X = 310 AND Y = 24 else
"000000000000" when X = 311 AND Y = 24 else
"000000000000" when X = 312 AND Y = 24 else
"000000000000" when X = 313 AND Y = 24 else
"000000000000" when X = 314 AND Y = 24 else
"000000000000" when X = 315 AND Y = 24 else
"000000000000" when X = 316 AND Y = 24 else
"000000000000" when X = 317 AND Y = 24 else
"000000000000" when X = 318 AND Y = 24 else
"000000000000" when X = 319 AND Y = 24 else
"000000000000" when X = 320 AND Y = 24 else
"000000000000" when X = 321 AND Y = 24 else
"000000000000" when X = 322 AND Y = 24 else
"000000000000" when X = 323 AND Y = 24 else
"000000000000" when X = 324 AND Y = 24 else
"000000000000" when X = 0 AND Y = 25 else
"000000000000" when X = 1 AND Y = 25 else
"000000000000" when X = 2 AND Y = 25 else
"000000000000" when X = 3 AND Y = 25 else
"000000000000" when X = 4 AND Y = 25 else
"000000000000" when X = 5 AND Y = 25 else
"000000000000" when X = 6 AND Y = 25 else
"000000000000" when X = 7 AND Y = 25 else
"000000000000" when X = 8 AND Y = 25 else
"000000000000" when X = 9 AND Y = 25 else
"000000000000" when X = 10 AND Y = 25 else
"000000000000" when X = 11 AND Y = 25 else
"000000000000" when X = 12 AND Y = 25 else
"000000000000" when X = 13 AND Y = 25 else
"000000000000" when X = 14 AND Y = 25 else
"000000000000" when X = 15 AND Y = 25 else
"000000000000" when X = 16 AND Y = 25 else
"000000000000" when X = 17 AND Y = 25 else
"000000000000" when X = 18 AND Y = 25 else
"000000000000" when X = 19 AND Y = 25 else
"000000000000" when X = 20 AND Y = 25 else
"000000000000" when X = 21 AND Y = 25 else
"000000000000" when X = 22 AND Y = 25 else
"000000000000" when X = 23 AND Y = 25 else
"000000000000" when X = 24 AND Y = 25 else
"000000000000" when X = 25 AND Y = 25 else
"000000000000" when X = 26 AND Y = 25 else
"000000000000" when X = 27 AND Y = 25 else
"000000000000" when X = 28 AND Y = 25 else
"000000000000" when X = 29 AND Y = 25 else
"000000000000" when X = 30 AND Y = 25 else
"000000000000" when X = 31 AND Y = 25 else
"000000000000" when X = 32 AND Y = 25 else
"000000000000" when X = 33 AND Y = 25 else
"000000000000" when X = 34 AND Y = 25 else
"000000000000" when X = 35 AND Y = 25 else
"000000000000" when X = 36 AND Y = 25 else
"000000000000" when X = 37 AND Y = 25 else
"000000000000" when X = 38 AND Y = 25 else
"000000000000" when X = 39 AND Y = 25 else
"100010011101" when X = 40 AND Y = 25 else
"100010011101" when X = 41 AND Y = 25 else
"100010011101" when X = 42 AND Y = 25 else
"100010011101" when X = 43 AND Y = 25 else
"100010011101" when X = 44 AND Y = 25 else
"100010011101" when X = 45 AND Y = 25 else
"100010011101" when X = 46 AND Y = 25 else
"100010011101" when X = 47 AND Y = 25 else
"100010011101" when X = 48 AND Y = 25 else
"100010011101" when X = 49 AND Y = 25 else
"110111011111" when X = 50 AND Y = 25 else
"110111011111" when X = 51 AND Y = 25 else
"110111011111" when X = 52 AND Y = 25 else
"110111011111" when X = 53 AND Y = 25 else
"110111011111" when X = 54 AND Y = 25 else
"110111011111" when X = 55 AND Y = 25 else
"110111011111" when X = 56 AND Y = 25 else
"110111011111" when X = 57 AND Y = 25 else
"110111011111" when X = 58 AND Y = 25 else
"110111011111" when X = 59 AND Y = 25 else
"111111111111" when X = 60 AND Y = 25 else
"111111111111" when X = 61 AND Y = 25 else
"111111111111" when X = 62 AND Y = 25 else
"111111111111" when X = 63 AND Y = 25 else
"111111111111" when X = 64 AND Y = 25 else
"111111111111" when X = 65 AND Y = 25 else
"111111111111" when X = 66 AND Y = 25 else
"111111111111" when X = 67 AND Y = 25 else
"111111111111" when X = 68 AND Y = 25 else
"111111111111" when X = 69 AND Y = 25 else
"111111111111" when X = 70 AND Y = 25 else
"111111111111" when X = 71 AND Y = 25 else
"111111111111" when X = 72 AND Y = 25 else
"111111111111" when X = 73 AND Y = 25 else
"111111111111" when X = 74 AND Y = 25 else
"111111111111" when X = 75 AND Y = 25 else
"111111111111" when X = 76 AND Y = 25 else
"111111111111" when X = 77 AND Y = 25 else
"111111111111" when X = 78 AND Y = 25 else
"111111111111" when X = 79 AND Y = 25 else
"111111111111" when X = 80 AND Y = 25 else
"111111111111" when X = 81 AND Y = 25 else
"111111111111" when X = 82 AND Y = 25 else
"111111111111" when X = 83 AND Y = 25 else
"111111111111" when X = 84 AND Y = 25 else
"111111111111" when X = 85 AND Y = 25 else
"111111111111" when X = 86 AND Y = 25 else
"111111111111" when X = 87 AND Y = 25 else
"111111111111" when X = 88 AND Y = 25 else
"111111111111" when X = 89 AND Y = 25 else
"111111111111" when X = 90 AND Y = 25 else
"111111111111" when X = 91 AND Y = 25 else
"111111111111" when X = 92 AND Y = 25 else
"111111111111" when X = 93 AND Y = 25 else
"111111111111" when X = 94 AND Y = 25 else
"111111111111" when X = 95 AND Y = 25 else
"111111111111" when X = 96 AND Y = 25 else
"111111111111" when X = 97 AND Y = 25 else
"111111111111" when X = 98 AND Y = 25 else
"111111111111" when X = 99 AND Y = 25 else
"111111111111" when X = 100 AND Y = 25 else
"111111111111" when X = 101 AND Y = 25 else
"111111111111" when X = 102 AND Y = 25 else
"111111111111" when X = 103 AND Y = 25 else
"111111111111" when X = 104 AND Y = 25 else
"111111111111" when X = 105 AND Y = 25 else
"111111111111" when X = 106 AND Y = 25 else
"111111111111" when X = 107 AND Y = 25 else
"111111111111" when X = 108 AND Y = 25 else
"111111111111" when X = 109 AND Y = 25 else
"111111111111" when X = 110 AND Y = 25 else
"111111111111" when X = 111 AND Y = 25 else
"111111111111" when X = 112 AND Y = 25 else
"111111111111" when X = 113 AND Y = 25 else
"111111111111" when X = 114 AND Y = 25 else
"111111111111" when X = 115 AND Y = 25 else
"111111111111" when X = 116 AND Y = 25 else
"111111111111" when X = 117 AND Y = 25 else
"111111111111" when X = 118 AND Y = 25 else
"111111111111" when X = 119 AND Y = 25 else
"111111111111" when X = 120 AND Y = 25 else
"111111111111" when X = 121 AND Y = 25 else
"111111111111" when X = 122 AND Y = 25 else
"111111111111" when X = 123 AND Y = 25 else
"111111111111" when X = 124 AND Y = 25 else
"111111111111" when X = 125 AND Y = 25 else
"111111111111" when X = 126 AND Y = 25 else
"111111111111" when X = 127 AND Y = 25 else
"111111111111" when X = 128 AND Y = 25 else
"111111111111" when X = 129 AND Y = 25 else
"111111111111" when X = 130 AND Y = 25 else
"111111111111" when X = 131 AND Y = 25 else
"111111111111" when X = 132 AND Y = 25 else
"111111111111" when X = 133 AND Y = 25 else
"111111111111" when X = 134 AND Y = 25 else
"111111111111" when X = 135 AND Y = 25 else
"111111111111" when X = 136 AND Y = 25 else
"111111111111" when X = 137 AND Y = 25 else
"111111111111" when X = 138 AND Y = 25 else
"111111111111" when X = 139 AND Y = 25 else
"111111111111" when X = 140 AND Y = 25 else
"111111111111" when X = 141 AND Y = 25 else
"111111111111" when X = 142 AND Y = 25 else
"111111111111" when X = 143 AND Y = 25 else
"111111111111" when X = 144 AND Y = 25 else
"111111111111" when X = 145 AND Y = 25 else
"111111111111" when X = 146 AND Y = 25 else
"111111111111" when X = 147 AND Y = 25 else
"111111111111" when X = 148 AND Y = 25 else
"111111111111" when X = 149 AND Y = 25 else
"111111111111" when X = 150 AND Y = 25 else
"111111111111" when X = 151 AND Y = 25 else
"111111111111" when X = 152 AND Y = 25 else
"111111111111" when X = 153 AND Y = 25 else
"111111111111" when X = 154 AND Y = 25 else
"111111111111" when X = 155 AND Y = 25 else
"111111111111" when X = 156 AND Y = 25 else
"111111111111" when X = 157 AND Y = 25 else
"111111111111" when X = 158 AND Y = 25 else
"111111111111" when X = 159 AND Y = 25 else
"000000000000" when X = 160 AND Y = 25 else
"000000000000" when X = 161 AND Y = 25 else
"000000000000" when X = 162 AND Y = 25 else
"000000000000" when X = 163 AND Y = 25 else
"000000000000" when X = 164 AND Y = 25 else
"000000000000" when X = 165 AND Y = 25 else
"000000000000" when X = 166 AND Y = 25 else
"000000000000" when X = 167 AND Y = 25 else
"000000000000" when X = 168 AND Y = 25 else
"000000000000" when X = 169 AND Y = 25 else
"000000000000" when X = 170 AND Y = 25 else
"000000000000" when X = 171 AND Y = 25 else
"000000000000" when X = 172 AND Y = 25 else
"000000000000" when X = 173 AND Y = 25 else
"000000000000" when X = 174 AND Y = 25 else
"000000000000" when X = 175 AND Y = 25 else
"000000000000" when X = 176 AND Y = 25 else
"000000000000" when X = 177 AND Y = 25 else
"000000000000" when X = 178 AND Y = 25 else
"000000000000" when X = 179 AND Y = 25 else
"000000000000" when X = 180 AND Y = 25 else
"000000000000" when X = 181 AND Y = 25 else
"000000000000" when X = 182 AND Y = 25 else
"000000000000" when X = 183 AND Y = 25 else
"000000000000" when X = 184 AND Y = 25 else
"000000000000" when X = 185 AND Y = 25 else
"000000000000" when X = 186 AND Y = 25 else
"000000000000" when X = 187 AND Y = 25 else
"000000000000" when X = 188 AND Y = 25 else
"000000000000" when X = 189 AND Y = 25 else
"000000000000" when X = 190 AND Y = 25 else
"000000000000" when X = 191 AND Y = 25 else
"000000000000" when X = 192 AND Y = 25 else
"000000000000" when X = 193 AND Y = 25 else
"000000000000" when X = 194 AND Y = 25 else
"000000000000" when X = 195 AND Y = 25 else
"000000000000" when X = 196 AND Y = 25 else
"000000000000" when X = 197 AND Y = 25 else
"000000000000" when X = 198 AND Y = 25 else
"000000000000" when X = 199 AND Y = 25 else
"000000000000" when X = 200 AND Y = 25 else
"000000000000" when X = 201 AND Y = 25 else
"000000000000" when X = 202 AND Y = 25 else
"000000000000" when X = 203 AND Y = 25 else
"000000000000" when X = 204 AND Y = 25 else
"000000000000" when X = 205 AND Y = 25 else
"000000000000" when X = 206 AND Y = 25 else
"000000000000" when X = 207 AND Y = 25 else
"000000000000" when X = 208 AND Y = 25 else
"000000000000" when X = 209 AND Y = 25 else
"000000000000" when X = 210 AND Y = 25 else
"000000000000" when X = 211 AND Y = 25 else
"000000000000" when X = 212 AND Y = 25 else
"000000000000" when X = 213 AND Y = 25 else
"000000000000" when X = 214 AND Y = 25 else
"000000000000" when X = 215 AND Y = 25 else
"000000000000" when X = 216 AND Y = 25 else
"000000000000" when X = 217 AND Y = 25 else
"000000000000" when X = 218 AND Y = 25 else
"000000000000" when X = 219 AND Y = 25 else
"000000000000" when X = 220 AND Y = 25 else
"000000000000" when X = 221 AND Y = 25 else
"000000000000" when X = 222 AND Y = 25 else
"000000000000" when X = 223 AND Y = 25 else
"000000000000" when X = 224 AND Y = 25 else
"000000000000" when X = 225 AND Y = 25 else
"000000000000" when X = 226 AND Y = 25 else
"000000000000" when X = 227 AND Y = 25 else
"000000000000" when X = 228 AND Y = 25 else
"000000000000" when X = 229 AND Y = 25 else
"000000000000" when X = 230 AND Y = 25 else
"000000000000" when X = 231 AND Y = 25 else
"000000000000" when X = 232 AND Y = 25 else
"000000000000" when X = 233 AND Y = 25 else
"000000000000" when X = 234 AND Y = 25 else
"111111111111" when X = 235 AND Y = 25 else
"111111111111" when X = 236 AND Y = 25 else
"111111111111" when X = 237 AND Y = 25 else
"111111111111" when X = 238 AND Y = 25 else
"111111111111" when X = 239 AND Y = 25 else
"111111111111" when X = 240 AND Y = 25 else
"111111111111" when X = 241 AND Y = 25 else
"111111111111" when X = 242 AND Y = 25 else
"111111111111" when X = 243 AND Y = 25 else
"111111111111" when X = 244 AND Y = 25 else
"111111111111" when X = 245 AND Y = 25 else
"111111111111" when X = 246 AND Y = 25 else
"111111111111" when X = 247 AND Y = 25 else
"111111111111" when X = 248 AND Y = 25 else
"111111111111" when X = 249 AND Y = 25 else
"110111011111" when X = 250 AND Y = 25 else
"110111011111" when X = 251 AND Y = 25 else
"110111011111" when X = 252 AND Y = 25 else
"110111011111" when X = 253 AND Y = 25 else
"110111011111" when X = 254 AND Y = 25 else
"110111011111" when X = 255 AND Y = 25 else
"110111011111" when X = 256 AND Y = 25 else
"110111011111" when X = 257 AND Y = 25 else
"110111011111" when X = 258 AND Y = 25 else
"110111011111" when X = 259 AND Y = 25 else
"110111011111" when X = 260 AND Y = 25 else
"110111011111" when X = 261 AND Y = 25 else
"110111011111" when X = 262 AND Y = 25 else
"110111011111" when X = 263 AND Y = 25 else
"110111011111" when X = 264 AND Y = 25 else
"110111011111" when X = 265 AND Y = 25 else
"110111011111" when X = 266 AND Y = 25 else
"110111011111" when X = 267 AND Y = 25 else
"110111011111" when X = 268 AND Y = 25 else
"110111011111" when X = 269 AND Y = 25 else
"110111011111" when X = 270 AND Y = 25 else
"110111011111" when X = 271 AND Y = 25 else
"110111011111" when X = 272 AND Y = 25 else
"110111011111" when X = 273 AND Y = 25 else
"110111011111" when X = 274 AND Y = 25 else
"110111011111" when X = 275 AND Y = 25 else
"110111011111" when X = 276 AND Y = 25 else
"110111011111" when X = 277 AND Y = 25 else
"110111011111" when X = 278 AND Y = 25 else
"110111011111" when X = 279 AND Y = 25 else
"000000000000" when X = 280 AND Y = 25 else
"000000000000" when X = 281 AND Y = 25 else
"000000000000" when X = 282 AND Y = 25 else
"000000000000" when X = 283 AND Y = 25 else
"000000000000" when X = 284 AND Y = 25 else
"000000000000" when X = 285 AND Y = 25 else
"000000000000" when X = 286 AND Y = 25 else
"000000000000" when X = 287 AND Y = 25 else
"000000000000" when X = 288 AND Y = 25 else
"000000000000" when X = 289 AND Y = 25 else
"000000000000" when X = 290 AND Y = 25 else
"000000000000" when X = 291 AND Y = 25 else
"000000000000" when X = 292 AND Y = 25 else
"000000000000" when X = 293 AND Y = 25 else
"000000000000" when X = 294 AND Y = 25 else
"000000000000" when X = 295 AND Y = 25 else
"000000000000" when X = 296 AND Y = 25 else
"000000000000" when X = 297 AND Y = 25 else
"000000000000" when X = 298 AND Y = 25 else
"000000000000" when X = 299 AND Y = 25 else
"000000000000" when X = 300 AND Y = 25 else
"000000000000" when X = 301 AND Y = 25 else
"000000000000" when X = 302 AND Y = 25 else
"000000000000" when X = 303 AND Y = 25 else
"000000000000" when X = 304 AND Y = 25 else
"000000000000" when X = 305 AND Y = 25 else
"000000000000" when X = 306 AND Y = 25 else
"000000000000" when X = 307 AND Y = 25 else
"000000000000" when X = 308 AND Y = 25 else
"000000000000" when X = 309 AND Y = 25 else
"000000000000" when X = 310 AND Y = 25 else
"000000000000" when X = 311 AND Y = 25 else
"000000000000" when X = 312 AND Y = 25 else
"000000000000" when X = 313 AND Y = 25 else
"000000000000" when X = 314 AND Y = 25 else
"000000000000" when X = 315 AND Y = 25 else
"000000000000" when X = 316 AND Y = 25 else
"000000000000" when X = 317 AND Y = 25 else
"000000000000" when X = 318 AND Y = 25 else
"000000000000" when X = 319 AND Y = 25 else
"000000000000" when X = 320 AND Y = 25 else
"000000000000" when X = 321 AND Y = 25 else
"000000000000" when X = 322 AND Y = 25 else
"000000000000" when X = 323 AND Y = 25 else
"000000000000" when X = 324 AND Y = 25 else
"000000000000" when X = 0 AND Y = 26 else
"000000000000" when X = 1 AND Y = 26 else
"000000000000" when X = 2 AND Y = 26 else
"000000000000" when X = 3 AND Y = 26 else
"000000000000" when X = 4 AND Y = 26 else
"000000000000" when X = 5 AND Y = 26 else
"000000000000" when X = 6 AND Y = 26 else
"000000000000" when X = 7 AND Y = 26 else
"000000000000" when X = 8 AND Y = 26 else
"000000000000" when X = 9 AND Y = 26 else
"000000000000" when X = 10 AND Y = 26 else
"000000000000" when X = 11 AND Y = 26 else
"000000000000" when X = 12 AND Y = 26 else
"000000000000" when X = 13 AND Y = 26 else
"000000000000" when X = 14 AND Y = 26 else
"000000000000" when X = 15 AND Y = 26 else
"000000000000" when X = 16 AND Y = 26 else
"000000000000" when X = 17 AND Y = 26 else
"000000000000" when X = 18 AND Y = 26 else
"000000000000" when X = 19 AND Y = 26 else
"000000000000" when X = 20 AND Y = 26 else
"000000000000" when X = 21 AND Y = 26 else
"000000000000" when X = 22 AND Y = 26 else
"000000000000" when X = 23 AND Y = 26 else
"000000000000" when X = 24 AND Y = 26 else
"000000000000" when X = 25 AND Y = 26 else
"000000000000" when X = 26 AND Y = 26 else
"000000000000" when X = 27 AND Y = 26 else
"000000000000" when X = 28 AND Y = 26 else
"000000000000" when X = 29 AND Y = 26 else
"000000000000" when X = 30 AND Y = 26 else
"000000000000" when X = 31 AND Y = 26 else
"000000000000" when X = 32 AND Y = 26 else
"000000000000" when X = 33 AND Y = 26 else
"000000000000" when X = 34 AND Y = 26 else
"000000000000" when X = 35 AND Y = 26 else
"000000000000" when X = 36 AND Y = 26 else
"000000000000" when X = 37 AND Y = 26 else
"000000000000" when X = 38 AND Y = 26 else
"000000000000" when X = 39 AND Y = 26 else
"100010011101" when X = 40 AND Y = 26 else
"100010011101" when X = 41 AND Y = 26 else
"100010011101" when X = 42 AND Y = 26 else
"100010011101" when X = 43 AND Y = 26 else
"100010011101" when X = 44 AND Y = 26 else
"100010011101" when X = 45 AND Y = 26 else
"100010011101" when X = 46 AND Y = 26 else
"100010011101" when X = 47 AND Y = 26 else
"100010011101" when X = 48 AND Y = 26 else
"100010011101" when X = 49 AND Y = 26 else
"110111011111" when X = 50 AND Y = 26 else
"110111011111" when X = 51 AND Y = 26 else
"110111011111" when X = 52 AND Y = 26 else
"110111011111" when X = 53 AND Y = 26 else
"110111011111" when X = 54 AND Y = 26 else
"110111011111" when X = 55 AND Y = 26 else
"110111011111" when X = 56 AND Y = 26 else
"110111011111" when X = 57 AND Y = 26 else
"110111011111" when X = 58 AND Y = 26 else
"110111011111" when X = 59 AND Y = 26 else
"111111111111" when X = 60 AND Y = 26 else
"111111111111" when X = 61 AND Y = 26 else
"111111111111" when X = 62 AND Y = 26 else
"111111111111" when X = 63 AND Y = 26 else
"111111111111" when X = 64 AND Y = 26 else
"111111111111" when X = 65 AND Y = 26 else
"111111111111" when X = 66 AND Y = 26 else
"111111111111" when X = 67 AND Y = 26 else
"111111111111" when X = 68 AND Y = 26 else
"111111111111" when X = 69 AND Y = 26 else
"111111111111" when X = 70 AND Y = 26 else
"111111111111" when X = 71 AND Y = 26 else
"111111111111" when X = 72 AND Y = 26 else
"111111111111" when X = 73 AND Y = 26 else
"111111111111" when X = 74 AND Y = 26 else
"111111111111" when X = 75 AND Y = 26 else
"111111111111" when X = 76 AND Y = 26 else
"111111111111" when X = 77 AND Y = 26 else
"111111111111" when X = 78 AND Y = 26 else
"111111111111" when X = 79 AND Y = 26 else
"111111111111" when X = 80 AND Y = 26 else
"111111111111" when X = 81 AND Y = 26 else
"111111111111" when X = 82 AND Y = 26 else
"111111111111" when X = 83 AND Y = 26 else
"111111111111" when X = 84 AND Y = 26 else
"111111111111" when X = 85 AND Y = 26 else
"111111111111" when X = 86 AND Y = 26 else
"111111111111" when X = 87 AND Y = 26 else
"111111111111" when X = 88 AND Y = 26 else
"111111111111" when X = 89 AND Y = 26 else
"111111111111" when X = 90 AND Y = 26 else
"111111111111" when X = 91 AND Y = 26 else
"111111111111" when X = 92 AND Y = 26 else
"111111111111" when X = 93 AND Y = 26 else
"111111111111" when X = 94 AND Y = 26 else
"111111111111" when X = 95 AND Y = 26 else
"111111111111" when X = 96 AND Y = 26 else
"111111111111" when X = 97 AND Y = 26 else
"111111111111" when X = 98 AND Y = 26 else
"111111111111" when X = 99 AND Y = 26 else
"111111111111" when X = 100 AND Y = 26 else
"111111111111" when X = 101 AND Y = 26 else
"111111111111" when X = 102 AND Y = 26 else
"111111111111" when X = 103 AND Y = 26 else
"111111111111" when X = 104 AND Y = 26 else
"111111111111" when X = 105 AND Y = 26 else
"111111111111" when X = 106 AND Y = 26 else
"111111111111" when X = 107 AND Y = 26 else
"111111111111" when X = 108 AND Y = 26 else
"111111111111" when X = 109 AND Y = 26 else
"111111111111" when X = 110 AND Y = 26 else
"111111111111" when X = 111 AND Y = 26 else
"111111111111" when X = 112 AND Y = 26 else
"111111111111" when X = 113 AND Y = 26 else
"111111111111" when X = 114 AND Y = 26 else
"111111111111" when X = 115 AND Y = 26 else
"111111111111" when X = 116 AND Y = 26 else
"111111111111" when X = 117 AND Y = 26 else
"111111111111" when X = 118 AND Y = 26 else
"111111111111" when X = 119 AND Y = 26 else
"111111111111" when X = 120 AND Y = 26 else
"111111111111" when X = 121 AND Y = 26 else
"111111111111" when X = 122 AND Y = 26 else
"111111111111" when X = 123 AND Y = 26 else
"111111111111" when X = 124 AND Y = 26 else
"111111111111" when X = 125 AND Y = 26 else
"111111111111" when X = 126 AND Y = 26 else
"111111111111" when X = 127 AND Y = 26 else
"111111111111" when X = 128 AND Y = 26 else
"111111111111" when X = 129 AND Y = 26 else
"111111111111" when X = 130 AND Y = 26 else
"111111111111" when X = 131 AND Y = 26 else
"111111111111" when X = 132 AND Y = 26 else
"111111111111" when X = 133 AND Y = 26 else
"111111111111" when X = 134 AND Y = 26 else
"111111111111" when X = 135 AND Y = 26 else
"111111111111" when X = 136 AND Y = 26 else
"111111111111" when X = 137 AND Y = 26 else
"111111111111" when X = 138 AND Y = 26 else
"111111111111" when X = 139 AND Y = 26 else
"111111111111" when X = 140 AND Y = 26 else
"111111111111" when X = 141 AND Y = 26 else
"111111111111" when X = 142 AND Y = 26 else
"111111111111" when X = 143 AND Y = 26 else
"111111111111" when X = 144 AND Y = 26 else
"111111111111" when X = 145 AND Y = 26 else
"111111111111" when X = 146 AND Y = 26 else
"111111111111" when X = 147 AND Y = 26 else
"111111111111" when X = 148 AND Y = 26 else
"111111111111" when X = 149 AND Y = 26 else
"111111111111" when X = 150 AND Y = 26 else
"111111111111" when X = 151 AND Y = 26 else
"111111111111" when X = 152 AND Y = 26 else
"111111111111" when X = 153 AND Y = 26 else
"111111111111" when X = 154 AND Y = 26 else
"111111111111" when X = 155 AND Y = 26 else
"111111111111" when X = 156 AND Y = 26 else
"111111111111" when X = 157 AND Y = 26 else
"111111111111" when X = 158 AND Y = 26 else
"111111111111" when X = 159 AND Y = 26 else
"000000000000" when X = 160 AND Y = 26 else
"000000000000" when X = 161 AND Y = 26 else
"000000000000" when X = 162 AND Y = 26 else
"000000000000" when X = 163 AND Y = 26 else
"000000000000" when X = 164 AND Y = 26 else
"000000000000" when X = 165 AND Y = 26 else
"000000000000" when X = 166 AND Y = 26 else
"000000000000" when X = 167 AND Y = 26 else
"000000000000" when X = 168 AND Y = 26 else
"000000000000" when X = 169 AND Y = 26 else
"000000000000" when X = 170 AND Y = 26 else
"000000000000" when X = 171 AND Y = 26 else
"000000000000" when X = 172 AND Y = 26 else
"000000000000" when X = 173 AND Y = 26 else
"000000000000" when X = 174 AND Y = 26 else
"000000000000" when X = 175 AND Y = 26 else
"000000000000" when X = 176 AND Y = 26 else
"000000000000" when X = 177 AND Y = 26 else
"000000000000" when X = 178 AND Y = 26 else
"000000000000" when X = 179 AND Y = 26 else
"000000000000" when X = 180 AND Y = 26 else
"000000000000" when X = 181 AND Y = 26 else
"000000000000" when X = 182 AND Y = 26 else
"000000000000" when X = 183 AND Y = 26 else
"000000000000" when X = 184 AND Y = 26 else
"000000000000" when X = 185 AND Y = 26 else
"000000000000" when X = 186 AND Y = 26 else
"000000000000" when X = 187 AND Y = 26 else
"000000000000" when X = 188 AND Y = 26 else
"000000000000" when X = 189 AND Y = 26 else
"000000000000" when X = 190 AND Y = 26 else
"000000000000" when X = 191 AND Y = 26 else
"000000000000" when X = 192 AND Y = 26 else
"000000000000" when X = 193 AND Y = 26 else
"000000000000" when X = 194 AND Y = 26 else
"000000000000" when X = 195 AND Y = 26 else
"000000000000" when X = 196 AND Y = 26 else
"000000000000" when X = 197 AND Y = 26 else
"000000000000" when X = 198 AND Y = 26 else
"000000000000" when X = 199 AND Y = 26 else
"000000000000" when X = 200 AND Y = 26 else
"000000000000" when X = 201 AND Y = 26 else
"000000000000" when X = 202 AND Y = 26 else
"000000000000" when X = 203 AND Y = 26 else
"000000000000" when X = 204 AND Y = 26 else
"000000000000" when X = 205 AND Y = 26 else
"000000000000" when X = 206 AND Y = 26 else
"000000000000" when X = 207 AND Y = 26 else
"000000000000" when X = 208 AND Y = 26 else
"000000000000" when X = 209 AND Y = 26 else
"000000000000" when X = 210 AND Y = 26 else
"000000000000" when X = 211 AND Y = 26 else
"000000000000" when X = 212 AND Y = 26 else
"000000000000" when X = 213 AND Y = 26 else
"000000000000" when X = 214 AND Y = 26 else
"000000000000" when X = 215 AND Y = 26 else
"000000000000" when X = 216 AND Y = 26 else
"000000000000" when X = 217 AND Y = 26 else
"000000000000" when X = 218 AND Y = 26 else
"000000000000" when X = 219 AND Y = 26 else
"000000000000" when X = 220 AND Y = 26 else
"000000000000" when X = 221 AND Y = 26 else
"000000000000" when X = 222 AND Y = 26 else
"000000000000" when X = 223 AND Y = 26 else
"000000000000" when X = 224 AND Y = 26 else
"000000000000" when X = 225 AND Y = 26 else
"000000000000" when X = 226 AND Y = 26 else
"000000000000" when X = 227 AND Y = 26 else
"000000000000" when X = 228 AND Y = 26 else
"000000000000" when X = 229 AND Y = 26 else
"000000000000" when X = 230 AND Y = 26 else
"000000000000" when X = 231 AND Y = 26 else
"000000000000" when X = 232 AND Y = 26 else
"000000000000" when X = 233 AND Y = 26 else
"000000000000" when X = 234 AND Y = 26 else
"111111111111" when X = 235 AND Y = 26 else
"111111111111" when X = 236 AND Y = 26 else
"111111111111" when X = 237 AND Y = 26 else
"111111111111" when X = 238 AND Y = 26 else
"111111111111" when X = 239 AND Y = 26 else
"111111111111" when X = 240 AND Y = 26 else
"111111111111" when X = 241 AND Y = 26 else
"111111111111" when X = 242 AND Y = 26 else
"111111111111" when X = 243 AND Y = 26 else
"111111111111" when X = 244 AND Y = 26 else
"111111111111" when X = 245 AND Y = 26 else
"111111111111" when X = 246 AND Y = 26 else
"111111111111" when X = 247 AND Y = 26 else
"111111111111" when X = 248 AND Y = 26 else
"111111111111" when X = 249 AND Y = 26 else
"110111011111" when X = 250 AND Y = 26 else
"110111011111" when X = 251 AND Y = 26 else
"110111011111" when X = 252 AND Y = 26 else
"110111011111" when X = 253 AND Y = 26 else
"110111011111" when X = 254 AND Y = 26 else
"110111011111" when X = 255 AND Y = 26 else
"110111011111" when X = 256 AND Y = 26 else
"110111011111" when X = 257 AND Y = 26 else
"110111011111" when X = 258 AND Y = 26 else
"110111011111" when X = 259 AND Y = 26 else
"110111011111" when X = 260 AND Y = 26 else
"110111011111" when X = 261 AND Y = 26 else
"110111011111" when X = 262 AND Y = 26 else
"110111011111" when X = 263 AND Y = 26 else
"110111011111" when X = 264 AND Y = 26 else
"110111011111" when X = 265 AND Y = 26 else
"110111011111" when X = 266 AND Y = 26 else
"110111011111" when X = 267 AND Y = 26 else
"110111011111" when X = 268 AND Y = 26 else
"110111011111" when X = 269 AND Y = 26 else
"110111011111" when X = 270 AND Y = 26 else
"110111011111" when X = 271 AND Y = 26 else
"110111011111" when X = 272 AND Y = 26 else
"110111011111" when X = 273 AND Y = 26 else
"110111011111" when X = 274 AND Y = 26 else
"110111011111" when X = 275 AND Y = 26 else
"110111011111" when X = 276 AND Y = 26 else
"110111011111" when X = 277 AND Y = 26 else
"110111011111" when X = 278 AND Y = 26 else
"110111011111" when X = 279 AND Y = 26 else
"000000000000" when X = 280 AND Y = 26 else
"000000000000" when X = 281 AND Y = 26 else
"000000000000" when X = 282 AND Y = 26 else
"000000000000" when X = 283 AND Y = 26 else
"000000000000" when X = 284 AND Y = 26 else
"000000000000" when X = 285 AND Y = 26 else
"000000000000" when X = 286 AND Y = 26 else
"000000000000" when X = 287 AND Y = 26 else
"000000000000" when X = 288 AND Y = 26 else
"000000000000" when X = 289 AND Y = 26 else
"000000000000" when X = 290 AND Y = 26 else
"000000000000" when X = 291 AND Y = 26 else
"000000000000" when X = 292 AND Y = 26 else
"000000000000" when X = 293 AND Y = 26 else
"000000000000" when X = 294 AND Y = 26 else
"000000000000" when X = 295 AND Y = 26 else
"000000000000" when X = 296 AND Y = 26 else
"000000000000" when X = 297 AND Y = 26 else
"000000000000" when X = 298 AND Y = 26 else
"000000000000" when X = 299 AND Y = 26 else
"000000000000" when X = 300 AND Y = 26 else
"000000000000" when X = 301 AND Y = 26 else
"000000000000" when X = 302 AND Y = 26 else
"000000000000" when X = 303 AND Y = 26 else
"000000000000" when X = 304 AND Y = 26 else
"000000000000" when X = 305 AND Y = 26 else
"000000000000" when X = 306 AND Y = 26 else
"000000000000" when X = 307 AND Y = 26 else
"000000000000" when X = 308 AND Y = 26 else
"000000000000" when X = 309 AND Y = 26 else
"000000000000" when X = 310 AND Y = 26 else
"000000000000" when X = 311 AND Y = 26 else
"000000000000" when X = 312 AND Y = 26 else
"000000000000" when X = 313 AND Y = 26 else
"000000000000" when X = 314 AND Y = 26 else
"000000000000" when X = 315 AND Y = 26 else
"000000000000" when X = 316 AND Y = 26 else
"000000000000" when X = 317 AND Y = 26 else
"000000000000" when X = 318 AND Y = 26 else
"000000000000" when X = 319 AND Y = 26 else
"000000000000" when X = 320 AND Y = 26 else
"000000000000" when X = 321 AND Y = 26 else
"000000000000" when X = 322 AND Y = 26 else
"000000000000" when X = 323 AND Y = 26 else
"000000000000" when X = 324 AND Y = 26 else
"000000000000" when X = 0 AND Y = 27 else
"000000000000" when X = 1 AND Y = 27 else
"000000000000" when X = 2 AND Y = 27 else
"000000000000" when X = 3 AND Y = 27 else
"000000000000" when X = 4 AND Y = 27 else
"000000000000" when X = 5 AND Y = 27 else
"000000000000" when X = 6 AND Y = 27 else
"000000000000" when X = 7 AND Y = 27 else
"000000000000" when X = 8 AND Y = 27 else
"000000000000" when X = 9 AND Y = 27 else
"000000000000" when X = 10 AND Y = 27 else
"000000000000" when X = 11 AND Y = 27 else
"000000000000" when X = 12 AND Y = 27 else
"000000000000" when X = 13 AND Y = 27 else
"000000000000" when X = 14 AND Y = 27 else
"000000000000" when X = 15 AND Y = 27 else
"000000000000" when X = 16 AND Y = 27 else
"000000000000" when X = 17 AND Y = 27 else
"000000000000" when X = 18 AND Y = 27 else
"000000000000" when X = 19 AND Y = 27 else
"000000000000" when X = 20 AND Y = 27 else
"000000000000" when X = 21 AND Y = 27 else
"000000000000" when X = 22 AND Y = 27 else
"000000000000" when X = 23 AND Y = 27 else
"000000000000" when X = 24 AND Y = 27 else
"000000000000" when X = 25 AND Y = 27 else
"000000000000" when X = 26 AND Y = 27 else
"000000000000" when X = 27 AND Y = 27 else
"000000000000" when X = 28 AND Y = 27 else
"000000000000" when X = 29 AND Y = 27 else
"000000000000" when X = 30 AND Y = 27 else
"000000000000" when X = 31 AND Y = 27 else
"000000000000" when X = 32 AND Y = 27 else
"000000000000" when X = 33 AND Y = 27 else
"000000000000" when X = 34 AND Y = 27 else
"000000000000" when X = 35 AND Y = 27 else
"000000000000" when X = 36 AND Y = 27 else
"000000000000" when X = 37 AND Y = 27 else
"000000000000" when X = 38 AND Y = 27 else
"000000000000" when X = 39 AND Y = 27 else
"100010011101" when X = 40 AND Y = 27 else
"100010011101" when X = 41 AND Y = 27 else
"100010011101" when X = 42 AND Y = 27 else
"100010011101" when X = 43 AND Y = 27 else
"100010011101" when X = 44 AND Y = 27 else
"100010011101" when X = 45 AND Y = 27 else
"100010011101" when X = 46 AND Y = 27 else
"100010011101" when X = 47 AND Y = 27 else
"100010011101" when X = 48 AND Y = 27 else
"100010011101" when X = 49 AND Y = 27 else
"110111011111" when X = 50 AND Y = 27 else
"110111011111" when X = 51 AND Y = 27 else
"110111011111" when X = 52 AND Y = 27 else
"110111011111" when X = 53 AND Y = 27 else
"110111011111" when X = 54 AND Y = 27 else
"110111011111" when X = 55 AND Y = 27 else
"110111011111" when X = 56 AND Y = 27 else
"110111011111" when X = 57 AND Y = 27 else
"110111011111" when X = 58 AND Y = 27 else
"110111011111" when X = 59 AND Y = 27 else
"111111111111" when X = 60 AND Y = 27 else
"111111111111" when X = 61 AND Y = 27 else
"111111111111" when X = 62 AND Y = 27 else
"111111111111" when X = 63 AND Y = 27 else
"111111111111" when X = 64 AND Y = 27 else
"111111111111" when X = 65 AND Y = 27 else
"111111111111" when X = 66 AND Y = 27 else
"111111111111" when X = 67 AND Y = 27 else
"111111111111" when X = 68 AND Y = 27 else
"111111111111" when X = 69 AND Y = 27 else
"111111111111" when X = 70 AND Y = 27 else
"111111111111" when X = 71 AND Y = 27 else
"111111111111" when X = 72 AND Y = 27 else
"111111111111" when X = 73 AND Y = 27 else
"111111111111" when X = 74 AND Y = 27 else
"111111111111" when X = 75 AND Y = 27 else
"111111111111" when X = 76 AND Y = 27 else
"111111111111" when X = 77 AND Y = 27 else
"111111111111" when X = 78 AND Y = 27 else
"111111111111" when X = 79 AND Y = 27 else
"111111111111" when X = 80 AND Y = 27 else
"111111111111" when X = 81 AND Y = 27 else
"111111111111" when X = 82 AND Y = 27 else
"111111111111" when X = 83 AND Y = 27 else
"111111111111" when X = 84 AND Y = 27 else
"111111111111" when X = 85 AND Y = 27 else
"111111111111" when X = 86 AND Y = 27 else
"111111111111" when X = 87 AND Y = 27 else
"111111111111" when X = 88 AND Y = 27 else
"111111111111" when X = 89 AND Y = 27 else
"111111111111" when X = 90 AND Y = 27 else
"111111111111" when X = 91 AND Y = 27 else
"111111111111" when X = 92 AND Y = 27 else
"111111111111" when X = 93 AND Y = 27 else
"111111111111" when X = 94 AND Y = 27 else
"111111111111" when X = 95 AND Y = 27 else
"111111111111" when X = 96 AND Y = 27 else
"111111111111" when X = 97 AND Y = 27 else
"111111111111" when X = 98 AND Y = 27 else
"111111111111" when X = 99 AND Y = 27 else
"111111111111" when X = 100 AND Y = 27 else
"111111111111" when X = 101 AND Y = 27 else
"111111111111" when X = 102 AND Y = 27 else
"111111111111" when X = 103 AND Y = 27 else
"111111111111" when X = 104 AND Y = 27 else
"111111111111" when X = 105 AND Y = 27 else
"111111111111" when X = 106 AND Y = 27 else
"111111111111" when X = 107 AND Y = 27 else
"111111111111" when X = 108 AND Y = 27 else
"111111111111" when X = 109 AND Y = 27 else
"111111111111" when X = 110 AND Y = 27 else
"111111111111" when X = 111 AND Y = 27 else
"111111111111" when X = 112 AND Y = 27 else
"111111111111" when X = 113 AND Y = 27 else
"111111111111" when X = 114 AND Y = 27 else
"111111111111" when X = 115 AND Y = 27 else
"111111111111" when X = 116 AND Y = 27 else
"111111111111" when X = 117 AND Y = 27 else
"111111111111" when X = 118 AND Y = 27 else
"111111111111" when X = 119 AND Y = 27 else
"111111111111" when X = 120 AND Y = 27 else
"111111111111" when X = 121 AND Y = 27 else
"111111111111" when X = 122 AND Y = 27 else
"111111111111" when X = 123 AND Y = 27 else
"111111111111" when X = 124 AND Y = 27 else
"111111111111" when X = 125 AND Y = 27 else
"111111111111" when X = 126 AND Y = 27 else
"111111111111" when X = 127 AND Y = 27 else
"111111111111" when X = 128 AND Y = 27 else
"111111111111" when X = 129 AND Y = 27 else
"111111111111" when X = 130 AND Y = 27 else
"111111111111" when X = 131 AND Y = 27 else
"111111111111" when X = 132 AND Y = 27 else
"111111111111" when X = 133 AND Y = 27 else
"111111111111" when X = 134 AND Y = 27 else
"111111111111" when X = 135 AND Y = 27 else
"111111111111" when X = 136 AND Y = 27 else
"111111111111" when X = 137 AND Y = 27 else
"111111111111" when X = 138 AND Y = 27 else
"111111111111" when X = 139 AND Y = 27 else
"111111111111" when X = 140 AND Y = 27 else
"111111111111" when X = 141 AND Y = 27 else
"111111111111" when X = 142 AND Y = 27 else
"111111111111" when X = 143 AND Y = 27 else
"111111111111" when X = 144 AND Y = 27 else
"111111111111" when X = 145 AND Y = 27 else
"111111111111" when X = 146 AND Y = 27 else
"111111111111" when X = 147 AND Y = 27 else
"111111111111" when X = 148 AND Y = 27 else
"111111111111" when X = 149 AND Y = 27 else
"111111111111" when X = 150 AND Y = 27 else
"111111111111" when X = 151 AND Y = 27 else
"111111111111" when X = 152 AND Y = 27 else
"111111111111" when X = 153 AND Y = 27 else
"111111111111" when X = 154 AND Y = 27 else
"111111111111" when X = 155 AND Y = 27 else
"111111111111" when X = 156 AND Y = 27 else
"111111111111" when X = 157 AND Y = 27 else
"111111111111" when X = 158 AND Y = 27 else
"111111111111" when X = 159 AND Y = 27 else
"000000000000" when X = 160 AND Y = 27 else
"000000000000" when X = 161 AND Y = 27 else
"000000000000" when X = 162 AND Y = 27 else
"000000000000" when X = 163 AND Y = 27 else
"000000000000" when X = 164 AND Y = 27 else
"000000000000" when X = 165 AND Y = 27 else
"000000000000" when X = 166 AND Y = 27 else
"000000000000" when X = 167 AND Y = 27 else
"000000000000" when X = 168 AND Y = 27 else
"000000000000" when X = 169 AND Y = 27 else
"000000000000" when X = 170 AND Y = 27 else
"000000000000" when X = 171 AND Y = 27 else
"000000000000" when X = 172 AND Y = 27 else
"000000000000" when X = 173 AND Y = 27 else
"000000000000" when X = 174 AND Y = 27 else
"000000000000" when X = 175 AND Y = 27 else
"000000000000" when X = 176 AND Y = 27 else
"000000000000" when X = 177 AND Y = 27 else
"000000000000" when X = 178 AND Y = 27 else
"000000000000" when X = 179 AND Y = 27 else
"000000000000" when X = 180 AND Y = 27 else
"000000000000" when X = 181 AND Y = 27 else
"000000000000" when X = 182 AND Y = 27 else
"000000000000" when X = 183 AND Y = 27 else
"000000000000" when X = 184 AND Y = 27 else
"000000000000" when X = 185 AND Y = 27 else
"000000000000" when X = 186 AND Y = 27 else
"000000000000" when X = 187 AND Y = 27 else
"000000000000" when X = 188 AND Y = 27 else
"000000000000" when X = 189 AND Y = 27 else
"000000000000" when X = 190 AND Y = 27 else
"000000000000" when X = 191 AND Y = 27 else
"000000000000" when X = 192 AND Y = 27 else
"000000000000" when X = 193 AND Y = 27 else
"000000000000" when X = 194 AND Y = 27 else
"000000000000" when X = 195 AND Y = 27 else
"000000000000" when X = 196 AND Y = 27 else
"000000000000" when X = 197 AND Y = 27 else
"000000000000" when X = 198 AND Y = 27 else
"000000000000" when X = 199 AND Y = 27 else
"000000000000" when X = 200 AND Y = 27 else
"000000000000" when X = 201 AND Y = 27 else
"000000000000" when X = 202 AND Y = 27 else
"000000000000" when X = 203 AND Y = 27 else
"000000000000" when X = 204 AND Y = 27 else
"000000000000" when X = 205 AND Y = 27 else
"000000000000" when X = 206 AND Y = 27 else
"000000000000" when X = 207 AND Y = 27 else
"000000000000" when X = 208 AND Y = 27 else
"000000000000" when X = 209 AND Y = 27 else
"000000000000" when X = 210 AND Y = 27 else
"000000000000" when X = 211 AND Y = 27 else
"000000000000" when X = 212 AND Y = 27 else
"000000000000" when X = 213 AND Y = 27 else
"000000000000" when X = 214 AND Y = 27 else
"000000000000" when X = 215 AND Y = 27 else
"000000000000" when X = 216 AND Y = 27 else
"000000000000" when X = 217 AND Y = 27 else
"000000000000" when X = 218 AND Y = 27 else
"000000000000" when X = 219 AND Y = 27 else
"000000000000" when X = 220 AND Y = 27 else
"000000000000" when X = 221 AND Y = 27 else
"000000000000" when X = 222 AND Y = 27 else
"000000000000" when X = 223 AND Y = 27 else
"000000000000" when X = 224 AND Y = 27 else
"000000000000" when X = 225 AND Y = 27 else
"000000000000" when X = 226 AND Y = 27 else
"000000000000" when X = 227 AND Y = 27 else
"000000000000" when X = 228 AND Y = 27 else
"000000000000" when X = 229 AND Y = 27 else
"000000000000" when X = 230 AND Y = 27 else
"000000000000" when X = 231 AND Y = 27 else
"000000000000" when X = 232 AND Y = 27 else
"000000000000" when X = 233 AND Y = 27 else
"000000000000" when X = 234 AND Y = 27 else
"111111111111" when X = 235 AND Y = 27 else
"111111111111" when X = 236 AND Y = 27 else
"111111111111" when X = 237 AND Y = 27 else
"111111111111" when X = 238 AND Y = 27 else
"111111111111" when X = 239 AND Y = 27 else
"111111111111" when X = 240 AND Y = 27 else
"111111111111" when X = 241 AND Y = 27 else
"111111111111" when X = 242 AND Y = 27 else
"111111111111" when X = 243 AND Y = 27 else
"111111111111" when X = 244 AND Y = 27 else
"111111111111" when X = 245 AND Y = 27 else
"111111111111" when X = 246 AND Y = 27 else
"111111111111" when X = 247 AND Y = 27 else
"111111111111" when X = 248 AND Y = 27 else
"111111111111" when X = 249 AND Y = 27 else
"110111011111" when X = 250 AND Y = 27 else
"110111011111" when X = 251 AND Y = 27 else
"110111011111" when X = 252 AND Y = 27 else
"110111011111" when X = 253 AND Y = 27 else
"110111011111" when X = 254 AND Y = 27 else
"110111011111" when X = 255 AND Y = 27 else
"110111011111" when X = 256 AND Y = 27 else
"110111011111" when X = 257 AND Y = 27 else
"110111011111" when X = 258 AND Y = 27 else
"110111011111" when X = 259 AND Y = 27 else
"110111011111" when X = 260 AND Y = 27 else
"110111011111" when X = 261 AND Y = 27 else
"110111011111" when X = 262 AND Y = 27 else
"110111011111" when X = 263 AND Y = 27 else
"110111011111" when X = 264 AND Y = 27 else
"110111011111" when X = 265 AND Y = 27 else
"110111011111" when X = 266 AND Y = 27 else
"110111011111" when X = 267 AND Y = 27 else
"110111011111" when X = 268 AND Y = 27 else
"110111011111" when X = 269 AND Y = 27 else
"110111011111" when X = 270 AND Y = 27 else
"110111011111" when X = 271 AND Y = 27 else
"110111011111" when X = 272 AND Y = 27 else
"110111011111" when X = 273 AND Y = 27 else
"110111011111" when X = 274 AND Y = 27 else
"110111011111" when X = 275 AND Y = 27 else
"110111011111" when X = 276 AND Y = 27 else
"110111011111" when X = 277 AND Y = 27 else
"110111011111" when X = 278 AND Y = 27 else
"110111011111" when X = 279 AND Y = 27 else
"000000000000" when X = 280 AND Y = 27 else
"000000000000" when X = 281 AND Y = 27 else
"000000000000" when X = 282 AND Y = 27 else
"000000000000" when X = 283 AND Y = 27 else
"000000000000" when X = 284 AND Y = 27 else
"000000000000" when X = 285 AND Y = 27 else
"000000000000" when X = 286 AND Y = 27 else
"000000000000" when X = 287 AND Y = 27 else
"000000000000" when X = 288 AND Y = 27 else
"000000000000" when X = 289 AND Y = 27 else
"000000000000" when X = 290 AND Y = 27 else
"000000000000" when X = 291 AND Y = 27 else
"000000000000" when X = 292 AND Y = 27 else
"000000000000" when X = 293 AND Y = 27 else
"000000000000" when X = 294 AND Y = 27 else
"000000000000" when X = 295 AND Y = 27 else
"000000000000" when X = 296 AND Y = 27 else
"000000000000" when X = 297 AND Y = 27 else
"000000000000" when X = 298 AND Y = 27 else
"000000000000" when X = 299 AND Y = 27 else
"000000000000" when X = 300 AND Y = 27 else
"000000000000" when X = 301 AND Y = 27 else
"000000000000" when X = 302 AND Y = 27 else
"000000000000" when X = 303 AND Y = 27 else
"000000000000" when X = 304 AND Y = 27 else
"000000000000" when X = 305 AND Y = 27 else
"000000000000" when X = 306 AND Y = 27 else
"000000000000" when X = 307 AND Y = 27 else
"000000000000" when X = 308 AND Y = 27 else
"000000000000" when X = 309 AND Y = 27 else
"000000000000" when X = 310 AND Y = 27 else
"000000000000" when X = 311 AND Y = 27 else
"000000000000" when X = 312 AND Y = 27 else
"000000000000" when X = 313 AND Y = 27 else
"000000000000" when X = 314 AND Y = 27 else
"000000000000" when X = 315 AND Y = 27 else
"000000000000" when X = 316 AND Y = 27 else
"000000000000" when X = 317 AND Y = 27 else
"000000000000" when X = 318 AND Y = 27 else
"000000000000" when X = 319 AND Y = 27 else
"000000000000" when X = 320 AND Y = 27 else
"000000000000" when X = 321 AND Y = 27 else
"000000000000" when X = 322 AND Y = 27 else
"000000000000" when X = 323 AND Y = 27 else
"000000000000" when X = 324 AND Y = 27 else
"000000000000" when X = 0 AND Y = 28 else
"000000000000" when X = 1 AND Y = 28 else
"000000000000" when X = 2 AND Y = 28 else
"000000000000" when X = 3 AND Y = 28 else
"000000000000" when X = 4 AND Y = 28 else
"000000000000" when X = 5 AND Y = 28 else
"000000000000" when X = 6 AND Y = 28 else
"000000000000" when X = 7 AND Y = 28 else
"000000000000" when X = 8 AND Y = 28 else
"000000000000" when X = 9 AND Y = 28 else
"000000000000" when X = 10 AND Y = 28 else
"000000000000" when X = 11 AND Y = 28 else
"000000000000" when X = 12 AND Y = 28 else
"000000000000" when X = 13 AND Y = 28 else
"000000000000" when X = 14 AND Y = 28 else
"000000000000" when X = 15 AND Y = 28 else
"000000000000" when X = 16 AND Y = 28 else
"000000000000" when X = 17 AND Y = 28 else
"000000000000" when X = 18 AND Y = 28 else
"000000000000" when X = 19 AND Y = 28 else
"000000000000" when X = 20 AND Y = 28 else
"000000000000" when X = 21 AND Y = 28 else
"000000000000" when X = 22 AND Y = 28 else
"000000000000" when X = 23 AND Y = 28 else
"000000000000" when X = 24 AND Y = 28 else
"000000000000" when X = 25 AND Y = 28 else
"000000000000" when X = 26 AND Y = 28 else
"000000000000" when X = 27 AND Y = 28 else
"000000000000" when X = 28 AND Y = 28 else
"000000000000" when X = 29 AND Y = 28 else
"000000000000" when X = 30 AND Y = 28 else
"000000000000" when X = 31 AND Y = 28 else
"000000000000" when X = 32 AND Y = 28 else
"000000000000" when X = 33 AND Y = 28 else
"000000000000" when X = 34 AND Y = 28 else
"000000000000" when X = 35 AND Y = 28 else
"000000000000" when X = 36 AND Y = 28 else
"000000000000" when X = 37 AND Y = 28 else
"000000000000" when X = 38 AND Y = 28 else
"000000000000" when X = 39 AND Y = 28 else
"100010011101" when X = 40 AND Y = 28 else
"100010011101" when X = 41 AND Y = 28 else
"100010011101" when X = 42 AND Y = 28 else
"100010011101" when X = 43 AND Y = 28 else
"100010011101" when X = 44 AND Y = 28 else
"100010011101" when X = 45 AND Y = 28 else
"100010011101" when X = 46 AND Y = 28 else
"100010011101" when X = 47 AND Y = 28 else
"100010011101" when X = 48 AND Y = 28 else
"100010011101" when X = 49 AND Y = 28 else
"110111011111" when X = 50 AND Y = 28 else
"110111011111" when X = 51 AND Y = 28 else
"110111011111" when X = 52 AND Y = 28 else
"110111011111" when X = 53 AND Y = 28 else
"110111011111" when X = 54 AND Y = 28 else
"110111011111" when X = 55 AND Y = 28 else
"110111011111" when X = 56 AND Y = 28 else
"110111011111" when X = 57 AND Y = 28 else
"110111011111" when X = 58 AND Y = 28 else
"110111011111" when X = 59 AND Y = 28 else
"111111111111" when X = 60 AND Y = 28 else
"111111111111" when X = 61 AND Y = 28 else
"111111111111" when X = 62 AND Y = 28 else
"111111111111" when X = 63 AND Y = 28 else
"111111111111" when X = 64 AND Y = 28 else
"111111111111" when X = 65 AND Y = 28 else
"111111111111" when X = 66 AND Y = 28 else
"111111111111" when X = 67 AND Y = 28 else
"111111111111" when X = 68 AND Y = 28 else
"111111111111" when X = 69 AND Y = 28 else
"111111111111" when X = 70 AND Y = 28 else
"111111111111" when X = 71 AND Y = 28 else
"111111111111" when X = 72 AND Y = 28 else
"111111111111" when X = 73 AND Y = 28 else
"111111111111" when X = 74 AND Y = 28 else
"111111111111" when X = 75 AND Y = 28 else
"111111111111" when X = 76 AND Y = 28 else
"111111111111" when X = 77 AND Y = 28 else
"111111111111" when X = 78 AND Y = 28 else
"111111111111" when X = 79 AND Y = 28 else
"111111111111" when X = 80 AND Y = 28 else
"111111111111" when X = 81 AND Y = 28 else
"111111111111" when X = 82 AND Y = 28 else
"111111111111" when X = 83 AND Y = 28 else
"111111111111" when X = 84 AND Y = 28 else
"111111111111" when X = 85 AND Y = 28 else
"111111111111" when X = 86 AND Y = 28 else
"111111111111" when X = 87 AND Y = 28 else
"111111111111" when X = 88 AND Y = 28 else
"111111111111" when X = 89 AND Y = 28 else
"111111111111" when X = 90 AND Y = 28 else
"111111111111" when X = 91 AND Y = 28 else
"111111111111" when X = 92 AND Y = 28 else
"111111111111" when X = 93 AND Y = 28 else
"111111111111" when X = 94 AND Y = 28 else
"111111111111" when X = 95 AND Y = 28 else
"111111111111" when X = 96 AND Y = 28 else
"111111111111" when X = 97 AND Y = 28 else
"111111111111" when X = 98 AND Y = 28 else
"111111111111" when X = 99 AND Y = 28 else
"111111111111" when X = 100 AND Y = 28 else
"111111111111" when X = 101 AND Y = 28 else
"111111111111" when X = 102 AND Y = 28 else
"111111111111" when X = 103 AND Y = 28 else
"111111111111" when X = 104 AND Y = 28 else
"111111111111" when X = 105 AND Y = 28 else
"111111111111" when X = 106 AND Y = 28 else
"111111111111" when X = 107 AND Y = 28 else
"111111111111" when X = 108 AND Y = 28 else
"111111111111" when X = 109 AND Y = 28 else
"111111111111" when X = 110 AND Y = 28 else
"111111111111" when X = 111 AND Y = 28 else
"111111111111" when X = 112 AND Y = 28 else
"111111111111" when X = 113 AND Y = 28 else
"111111111111" when X = 114 AND Y = 28 else
"111111111111" when X = 115 AND Y = 28 else
"111111111111" when X = 116 AND Y = 28 else
"111111111111" when X = 117 AND Y = 28 else
"111111111111" when X = 118 AND Y = 28 else
"111111111111" when X = 119 AND Y = 28 else
"111111111111" when X = 120 AND Y = 28 else
"111111111111" when X = 121 AND Y = 28 else
"111111111111" when X = 122 AND Y = 28 else
"111111111111" when X = 123 AND Y = 28 else
"111111111111" when X = 124 AND Y = 28 else
"111111111111" when X = 125 AND Y = 28 else
"111111111111" when X = 126 AND Y = 28 else
"111111111111" when X = 127 AND Y = 28 else
"111111111111" when X = 128 AND Y = 28 else
"111111111111" when X = 129 AND Y = 28 else
"111111111111" when X = 130 AND Y = 28 else
"111111111111" when X = 131 AND Y = 28 else
"111111111111" when X = 132 AND Y = 28 else
"111111111111" when X = 133 AND Y = 28 else
"111111111111" when X = 134 AND Y = 28 else
"111111111111" when X = 135 AND Y = 28 else
"111111111111" when X = 136 AND Y = 28 else
"111111111111" when X = 137 AND Y = 28 else
"111111111111" when X = 138 AND Y = 28 else
"111111111111" when X = 139 AND Y = 28 else
"111111111111" when X = 140 AND Y = 28 else
"111111111111" when X = 141 AND Y = 28 else
"111111111111" when X = 142 AND Y = 28 else
"111111111111" when X = 143 AND Y = 28 else
"111111111111" when X = 144 AND Y = 28 else
"111111111111" when X = 145 AND Y = 28 else
"111111111111" when X = 146 AND Y = 28 else
"111111111111" when X = 147 AND Y = 28 else
"111111111111" when X = 148 AND Y = 28 else
"111111111111" when X = 149 AND Y = 28 else
"111111111111" when X = 150 AND Y = 28 else
"111111111111" when X = 151 AND Y = 28 else
"111111111111" when X = 152 AND Y = 28 else
"111111111111" when X = 153 AND Y = 28 else
"111111111111" when X = 154 AND Y = 28 else
"111111111111" when X = 155 AND Y = 28 else
"111111111111" when X = 156 AND Y = 28 else
"111111111111" when X = 157 AND Y = 28 else
"111111111111" when X = 158 AND Y = 28 else
"111111111111" when X = 159 AND Y = 28 else
"000000000000" when X = 160 AND Y = 28 else
"000000000000" when X = 161 AND Y = 28 else
"000000000000" when X = 162 AND Y = 28 else
"000000000000" when X = 163 AND Y = 28 else
"000000000000" when X = 164 AND Y = 28 else
"000000000000" when X = 165 AND Y = 28 else
"000000000000" when X = 166 AND Y = 28 else
"000000000000" when X = 167 AND Y = 28 else
"000000000000" when X = 168 AND Y = 28 else
"000000000000" when X = 169 AND Y = 28 else
"000000000000" when X = 170 AND Y = 28 else
"000000000000" when X = 171 AND Y = 28 else
"000000000000" when X = 172 AND Y = 28 else
"000000000000" when X = 173 AND Y = 28 else
"000000000000" when X = 174 AND Y = 28 else
"000000000000" when X = 175 AND Y = 28 else
"000000000000" when X = 176 AND Y = 28 else
"000000000000" when X = 177 AND Y = 28 else
"000000000000" when X = 178 AND Y = 28 else
"000000000000" when X = 179 AND Y = 28 else
"000000000000" when X = 180 AND Y = 28 else
"000000000000" when X = 181 AND Y = 28 else
"000000000000" when X = 182 AND Y = 28 else
"000000000000" when X = 183 AND Y = 28 else
"000000000000" when X = 184 AND Y = 28 else
"000000000000" when X = 185 AND Y = 28 else
"000000000000" when X = 186 AND Y = 28 else
"000000000000" when X = 187 AND Y = 28 else
"000000000000" when X = 188 AND Y = 28 else
"000000000000" when X = 189 AND Y = 28 else
"000000000000" when X = 190 AND Y = 28 else
"000000000000" when X = 191 AND Y = 28 else
"000000000000" when X = 192 AND Y = 28 else
"000000000000" when X = 193 AND Y = 28 else
"000000000000" when X = 194 AND Y = 28 else
"000000000000" when X = 195 AND Y = 28 else
"000000000000" when X = 196 AND Y = 28 else
"000000000000" when X = 197 AND Y = 28 else
"000000000000" when X = 198 AND Y = 28 else
"000000000000" when X = 199 AND Y = 28 else
"000000000000" when X = 200 AND Y = 28 else
"000000000000" when X = 201 AND Y = 28 else
"000000000000" when X = 202 AND Y = 28 else
"000000000000" when X = 203 AND Y = 28 else
"000000000000" when X = 204 AND Y = 28 else
"000000000000" when X = 205 AND Y = 28 else
"000000000000" when X = 206 AND Y = 28 else
"000000000000" when X = 207 AND Y = 28 else
"000000000000" when X = 208 AND Y = 28 else
"000000000000" when X = 209 AND Y = 28 else
"000000000000" when X = 210 AND Y = 28 else
"000000000000" when X = 211 AND Y = 28 else
"000000000000" when X = 212 AND Y = 28 else
"000000000000" when X = 213 AND Y = 28 else
"000000000000" when X = 214 AND Y = 28 else
"000000000000" when X = 215 AND Y = 28 else
"000000000000" when X = 216 AND Y = 28 else
"000000000000" when X = 217 AND Y = 28 else
"000000000000" when X = 218 AND Y = 28 else
"000000000000" when X = 219 AND Y = 28 else
"000000000000" when X = 220 AND Y = 28 else
"000000000000" when X = 221 AND Y = 28 else
"000000000000" when X = 222 AND Y = 28 else
"000000000000" when X = 223 AND Y = 28 else
"000000000000" when X = 224 AND Y = 28 else
"000000000000" when X = 225 AND Y = 28 else
"000000000000" when X = 226 AND Y = 28 else
"000000000000" when X = 227 AND Y = 28 else
"000000000000" when X = 228 AND Y = 28 else
"000000000000" when X = 229 AND Y = 28 else
"000000000000" when X = 230 AND Y = 28 else
"000000000000" when X = 231 AND Y = 28 else
"000000000000" when X = 232 AND Y = 28 else
"000000000000" when X = 233 AND Y = 28 else
"000000000000" when X = 234 AND Y = 28 else
"111111111111" when X = 235 AND Y = 28 else
"111111111111" when X = 236 AND Y = 28 else
"111111111111" when X = 237 AND Y = 28 else
"111111111111" when X = 238 AND Y = 28 else
"111111111111" when X = 239 AND Y = 28 else
"111111111111" when X = 240 AND Y = 28 else
"111111111111" when X = 241 AND Y = 28 else
"111111111111" when X = 242 AND Y = 28 else
"111111111111" when X = 243 AND Y = 28 else
"111111111111" when X = 244 AND Y = 28 else
"111111111111" when X = 245 AND Y = 28 else
"111111111111" when X = 246 AND Y = 28 else
"111111111111" when X = 247 AND Y = 28 else
"111111111111" when X = 248 AND Y = 28 else
"111111111111" when X = 249 AND Y = 28 else
"110111011111" when X = 250 AND Y = 28 else
"110111011111" when X = 251 AND Y = 28 else
"110111011111" when X = 252 AND Y = 28 else
"110111011111" when X = 253 AND Y = 28 else
"110111011111" when X = 254 AND Y = 28 else
"110111011111" when X = 255 AND Y = 28 else
"110111011111" when X = 256 AND Y = 28 else
"110111011111" when X = 257 AND Y = 28 else
"110111011111" when X = 258 AND Y = 28 else
"110111011111" when X = 259 AND Y = 28 else
"110111011111" when X = 260 AND Y = 28 else
"110111011111" when X = 261 AND Y = 28 else
"110111011111" when X = 262 AND Y = 28 else
"110111011111" when X = 263 AND Y = 28 else
"110111011111" when X = 264 AND Y = 28 else
"110111011111" when X = 265 AND Y = 28 else
"110111011111" when X = 266 AND Y = 28 else
"110111011111" when X = 267 AND Y = 28 else
"110111011111" when X = 268 AND Y = 28 else
"110111011111" when X = 269 AND Y = 28 else
"110111011111" when X = 270 AND Y = 28 else
"110111011111" when X = 271 AND Y = 28 else
"110111011111" when X = 272 AND Y = 28 else
"110111011111" when X = 273 AND Y = 28 else
"110111011111" when X = 274 AND Y = 28 else
"110111011111" when X = 275 AND Y = 28 else
"110111011111" when X = 276 AND Y = 28 else
"110111011111" when X = 277 AND Y = 28 else
"110111011111" when X = 278 AND Y = 28 else
"110111011111" when X = 279 AND Y = 28 else
"000000000000" when X = 280 AND Y = 28 else
"000000000000" when X = 281 AND Y = 28 else
"000000000000" when X = 282 AND Y = 28 else
"000000000000" when X = 283 AND Y = 28 else
"000000000000" when X = 284 AND Y = 28 else
"000000000000" when X = 285 AND Y = 28 else
"000000000000" when X = 286 AND Y = 28 else
"000000000000" when X = 287 AND Y = 28 else
"000000000000" when X = 288 AND Y = 28 else
"000000000000" when X = 289 AND Y = 28 else
"000000000000" when X = 290 AND Y = 28 else
"000000000000" when X = 291 AND Y = 28 else
"000000000000" when X = 292 AND Y = 28 else
"000000000000" when X = 293 AND Y = 28 else
"000000000000" when X = 294 AND Y = 28 else
"000000000000" when X = 295 AND Y = 28 else
"000000000000" when X = 296 AND Y = 28 else
"000000000000" when X = 297 AND Y = 28 else
"000000000000" when X = 298 AND Y = 28 else
"000000000000" when X = 299 AND Y = 28 else
"000000000000" when X = 300 AND Y = 28 else
"000000000000" when X = 301 AND Y = 28 else
"000000000000" when X = 302 AND Y = 28 else
"000000000000" when X = 303 AND Y = 28 else
"000000000000" when X = 304 AND Y = 28 else
"000000000000" when X = 305 AND Y = 28 else
"000000000000" when X = 306 AND Y = 28 else
"000000000000" when X = 307 AND Y = 28 else
"000000000000" when X = 308 AND Y = 28 else
"000000000000" when X = 309 AND Y = 28 else
"000000000000" when X = 310 AND Y = 28 else
"000000000000" when X = 311 AND Y = 28 else
"000000000000" when X = 312 AND Y = 28 else
"000000000000" when X = 313 AND Y = 28 else
"000000000000" when X = 314 AND Y = 28 else
"000000000000" when X = 315 AND Y = 28 else
"000000000000" when X = 316 AND Y = 28 else
"000000000000" when X = 317 AND Y = 28 else
"000000000000" when X = 318 AND Y = 28 else
"000000000000" when X = 319 AND Y = 28 else
"000000000000" when X = 320 AND Y = 28 else
"000000000000" when X = 321 AND Y = 28 else
"000000000000" when X = 322 AND Y = 28 else
"000000000000" when X = 323 AND Y = 28 else
"000000000000" when X = 324 AND Y = 28 else
"000000000000" when X = 0 AND Y = 29 else
"000000000000" when X = 1 AND Y = 29 else
"000000000000" when X = 2 AND Y = 29 else
"000000000000" when X = 3 AND Y = 29 else
"000000000000" when X = 4 AND Y = 29 else
"000000000000" when X = 5 AND Y = 29 else
"000000000000" when X = 6 AND Y = 29 else
"000000000000" when X = 7 AND Y = 29 else
"000000000000" when X = 8 AND Y = 29 else
"000000000000" when X = 9 AND Y = 29 else
"000000000000" when X = 10 AND Y = 29 else
"000000000000" when X = 11 AND Y = 29 else
"000000000000" when X = 12 AND Y = 29 else
"000000000000" when X = 13 AND Y = 29 else
"000000000000" when X = 14 AND Y = 29 else
"000000000000" when X = 15 AND Y = 29 else
"000000000000" when X = 16 AND Y = 29 else
"000000000000" when X = 17 AND Y = 29 else
"000000000000" when X = 18 AND Y = 29 else
"000000000000" when X = 19 AND Y = 29 else
"000000000000" when X = 20 AND Y = 29 else
"000000000000" when X = 21 AND Y = 29 else
"000000000000" when X = 22 AND Y = 29 else
"000000000000" when X = 23 AND Y = 29 else
"000000000000" when X = 24 AND Y = 29 else
"000000000000" when X = 25 AND Y = 29 else
"000000000000" when X = 26 AND Y = 29 else
"000000000000" when X = 27 AND Y = 29 else
"000000000000" when X = 28 AND Y = 29 else
"000000000000" when X = 29 AND Y = 29 else
"000000000000" when X = 30 AND Y = 29 else
"000000000000" when X = 31 AND Y = 29 else
"000000000000" when X = 32 AND Y = 29 else
"000000000000" when X = 33 AND Y = 29 else
"000000000000" when X = 34 AND Y = 29 else
"000000000000" when X = 35 AND Y = 29 else
"000000000000" when X = 36 AND Y = 29 else
"000000000000" when X = 37 AND Y = 29 else
"000000000000" when X = 38 AND Y = 29 else
"000000000000" when X = 39 AND Y = 29 else
"100010011101" when X = 40 AND Y = 29 else
"100010011101" when X = 41 AND Y = 29 else
"100010011101" when X = 42 AND Y = 29 else
"100010011101" when X = 43 AND Y = 29 else
"100010011101" when X = 44 AND Y = 29 else
"100010011101" when X = 45 AND Y = 29 else
"100010011101" when X = 46 AND Y = 29 else
"100010011101" when X = 47 AND Y = 29 else
"100010011101" when X = 48 AND Y = 29 else
"100010011101" when X = 49 AND Y = 29 else
"110111011111" when X = 50 AND Y = 29 else
"110111011111" when X = 51 AND Y = 29 else
"110111011111" when X = 52 AND Y = 29 else
"110111011111" when X = 53 AND Y = 29 else
"110111011111" when X = 54 AND Y = 29 else
"110111011111" when X = 55 AND Y = 29 else
"110111011111" when X = 56 AND Y = 29 else
"110111011111" when X = 57 AND Y = 29 else
"110111011111" when X = 58 AND Y = 29 else
"110111011111" when X = 59 AND Y = 29 else
"111111111111" when X = 60 AND Y = 29 else
"111111111111" when X = 61 AND Y = 29 else
"111111111111" when X = 62 AND Y = 29 else
"111111111111" when X = 63 AND Y = 29 else
"111111111111" when X = 64 AND Y = 29 else
"111111111111" when X = 65 AND Y = 29 else
"111111111111" when X = 66 AND Y = 29 else
"111111111111" when X = 67 AND Y = 29 else
"111111111111" when X = 68 AND Y = 29 else
"111111111111" when X = 69 AND Y = 29 else
"111111111111" when X = 70 AND Y = 29 else
"111111111111" when X = 71 AND Y = 29 else
"111111111111" when X = 72 AND Y = 29 else
"111111111111" when X = 73 AND Y = 29 else
"111111111111" when X = 74 AND Y = 29 else
"111111111111" when X = 75 AND Y = 29 else
"111111111111" when X = 76 AND Y = 29 else
"111111111111" when X = 77 AND Y = 29 else
"111111111111" when X = 78 AND Y = 29 else
"111111111111" when X = 79 AND Y = 29 else
"111111111111" when X = 80 AND Y = 29 else
"111111111111" when X = 81 AND Y = 29 else
"111111111111" when X = 82 AND Y = 29 else
"111111111111" when X = 83 AND Y = 29 else
"111111111111" when X = 84 AND Y = 29 else
"111111111111" when X = 85 AND Y = 29 else
"111111111111" when X = 86 AND Y = 29 else
"111111111111" when X = 87 AND Y = 29 else
"111111111111" when X = 88 AND Y = 29 else
"111111111111" when X = 89 AND Y = 29 else
"111111111111" when X = 90 AND Y = 29 else
"111111111111" when X = 91 AND Y = 29 else
"111111111111" when X = 92 AND Y = 29 else
"111111111111" when X = 93 AND Y = 29 else
"111111111111" when X = 94 AND Y = 29 else
"111111111111" when X = 95 AND Y = 29 else
"111111111111" when X = 96 AND Y = 29 else
"111111111111" when X = 97 AND Y = 29 else
"111111111111" when X = 98 AND Y = 29 else
"111111111111" when X = 99 AND Y = 29 else
"111111111111" when X = 100 AND Y = 29 else
"111111111111" when X = 101 AND Y = 29 else
"111111111111" when X = 102 AND Y = 29 else
"111111111111" when X = 103 AND Y = 29 else
"111111111111" when X = 104 AND Y = 29 else
"111111111111" when X = 105 AND Y = 29 else
"111111111111" when X = 106 AND Y = 29 else
"111111111111" when X = 107 AND Y = 29 else
"111111111111" when X = 108 AND Y = 29 else
"111111111111" when X = 109 AND Y = 29 else
"111111111111" when X = 110 AND Y = 29 else
"111111111111" when X = 111 AND Y = 29 else
"111111111111" when X = 112 AND Y = 29 else
"111111111111" when X = 113 AND Y = 29 else
"111111111111" when X = 114 AND Y = 29 else
"111111111111" when X = 115 AND Y = 29 else
"111111111111" when X = 116 AND Y = 29 else
"111111111111" when X = 117 AND Y = 29 else
"111111111111" when X = 118 AND Y = 29 else
"111111111111" when X = 119 AND Y = 29 else
"111111111111" when X = 120 AND Y = 29 else
"111111111111" when X = 121 AND Y = 29 else
"111111111111" when X = 122 AND Y = 29 else
"111111111111" when X = 123 AND Y = 29 else
"111111111111" when X = 124 AND Y = 29 else
"111111111111" when X = 125 AND Y = 29 else
"111111111111" when X = 126 AND Y = 29 else
"111111111111" when X = 127 AND Y = 29 else
"111111111111" when X = 128 AND Y = 29 else
"111111111111" when X = 129 AND Y = 29 else
"111111111111" when X = 130 AND Y = 29 else
"111111111111" when X = 131 AND Y = 29 else
"111111111111" when X = 132 AND Y = 29 else
"111111111111" when X = 133 AND Y = 29 else
"111111111111" when X = 134 AND Y = 29 else
"111111111111" when X = 135 AND Y = 29 else
"111111111111" when X = 136 AND Y = 29 else
"111111111111" when X = 137 AND Y = 29 else
"111111111111" when X = 138 AND Y = 29 else
"111111111111" when X = 139 AND Y = 29 else
"111111111111" when X = 140 AND Y = 29 else
"111111111111" when X = 141 AND Y = 29 else
"111111111111" when X = 142 AND Y = 29 else
"111111111111" when X = 143 AND Y = 29 else
"111111111111" when X = 144 AND Y = 29 else
"111111111111" when X = 145 AND Y = 29 else
"111111111111" when X = 146 AND Y = 29 else
"111111111111" when X = 147 AND Y = 29 else
"111111111111" when X = 148 AND Y = 29 else
"111111111111" when X = 149 AND Y = 29 else
"111111111111" when X = 150 AND Y = 29 else
"111111111111" when X = 151 AND Y = 29 else
"111111111111" when X = 152 AND Y = 29 else
"111111111111" when X = 153 AND Y = 29 else
"111111111111" when X = 154 AND Y = 29 else
"111111111111" when X = 155 AND Y = 29 else
"111111111111" when X = 156 AND Y = 29 else
"111111111111" when X = 157 AND Y = 29 else
"111111111111" when X = 158 AND Y = 29 else
"111111111111" when X = 159 AND Y = 29 else
"000000000000" when X = 160 AND Y = 29 else
"000000000000" when X = 161 AND Y = 29 else
"000000000000" when X = 162 AND Y = 29 else
"000000000000" when X = 163 AND Y = 29 else
"000000000000" when X = 164 AND Y = 29 else
"000000000000" when X = 165 AND Y = 29 else
"000000000000" when X = 166 AND Y = 29 else
"000000000000" when X = 167 AND Y = 29 else
"000000000000" when X = 168 AND Y = 29 else
"000000000000" when X = 169 AND Y = 29 else
"000000000000" when X = 170 AND Y = 29 else
"000000000000" when X = 171 AND Y = 29 else
"000000000000" when X = 172 AND Y = 29 else
"000000000000" when X = 173 AND Y = 29 else
"000000000000" when X = 174 AND Y = 29 else
"000000000000" when X = 175 AND Y = 29 else
"000000000000" when X = 176 AND Y = 29 else
"000000000000" when X = 177 AND Y = 29 else
"000000000000" when X = 178 AND Y = 29 else
"000000000000" when X = 179 AND Y = 29 else
"000000000000" when X = 180 AND Y = 29 else
"000000000000" when X = 181 AND Y = 29 else
"000000000000" when X = 182 AND Y = 29 else
"000000000000" when X = 183 AND Y = 29 else
"000000000000" when X = 184 AND Y = 29 else
"000000000000" when X = 185 AND Y = 29 else
"000000000000" when X = 186 AND Y = 29 else
"000000000000" when X = 187 AND Y = 29 else
"000000000000" when X = 188 AND Y = 29 else
"000000000000" when X = 189 AND Y = 29 else
"000000000000" when X = 190 AND Y = 29 else
"000000000000" when X = 191 AND Y = 29 else
"000000000000" when X = 192 AND Y = 29 else
"000000000000" when X = 193 AND Y = 29 else
"000000000000" when X = 194 AND Y = 29 else
"000000000000" when X = 195 AND Y = 29 else
"000000000000" when X = 196 AND Y = 29 else
"000000000000" when X = 197 AND Y = 29 else
"000000000000" when X = 198 AND Y = 29 else
"000000000000" when X = 199 AND Y = 29 else
"000000000000" when X = 200 AND Y = 29 else
"000000000000" when X = 201 AND Y = 29 else
"000000000000" when X = 202 AND Y = 29 else
"000000000000" when X = 203 AND Y = 29 else
"000000000000" when X = 204 AND Y = 29 else
"000000000000" when X = 205 AND Y = 29 else
"000000000000" when X = 206 AND Y = 29 else
"000000000000" when X = 207 AND Y = 29 else
"000000000000" when X = 208 AND Y = 29 else
"000000000000" when X = 209 AND Y = 29 else
"000000000000" when X = 210 AND Y = 29 else
"000000000000" when X = 211 AND Y = 29 else
"000000000000" when X = 212 AND Y = 29 else
"000000000000" when X = 213 AND Y = 29 else
"000000000000" when X = 214 AND Y = 29 else
"000000000000" when X = 215 AND Y = 29 else
"000000000000" when X = 216 AND Y = 29 else
"000000000000" when X = 217 AND Y = 29 else
"000000000000" when X = 218 AND Y = 29 else
"000000000000" when X = 219 AND Y = 29 else
"000000000000" when X = 220 AND Y = 29 else
"000000000000" when X = 221 AND Y = 29 else
"000000000000" when X = 222 AND Y = 29 else
"000000000000" when X = 223 AND Y = 29 else
"000000000000" when X = 224 AND Y = 29 else
"000000000000" when X = 225 AND Y = 29 else
"000000000000" when X = 226 AND Y = 29 else
"000000000000" when X = 227 AND Y = 29 else
"000000000000" when X = 228 AND Y = 29 else
"000000000000" when X = 229 AND Y = 29 else
"000000000000" when X = 230 AND Y = 29 else
"000000000000" when X = 231 AND Y = 29 else
"000000000000" when X = 232 AND Y = 29 else
"000000000000" when X = 233 AND Y = 29 else
"000000000000" when X = 234 AND Y = 29 else
"111111111111" when X = 235 AND Y = 29 else
"111111111111" when X = 236 AND Y = 29 else
"111111111111" when X = 237 AND Y = 29 else
"111111111111" when X = 238 AND Y = 29 else
"111111111111" when X = 239 AND Y = 29 else
"111111111111" when X = 240 AND Y = 29 else
"111111111111" when X = 241 AND Y = 29 else
"111111111111" when X = 242 AND Y = 29 else
"111111111111" when X = 243 AND Y = 29 else
"111111111111" when X = 244 AND Y = 29 else
"111111111111" when X = 245 AND Y = 29 else
"111111111111" when X = 246 AND Y = 29 else
"111111111111" when X = 247 AND Y = 29 else
"111111111111" when X = 248 AND Y = 29 else
"111111111111" when X = 249 AND Y = 29 else
"110111011111" when X = 250 AND Y = 29 else
"110111011111" when X = 251 AND Y = 29 else
"110111011111" when X = 252 AND Y = 29 else
"110111011111" when X = 253 AND Y = 29 else
"110111011111" when X = 254 AND Y = 29 else
"110111011111" when X = 255 AND Y = 29 else
"110111011111" when X = 256 AND Y = 29 else
"110111011111" when X = 257 AND Y = 29 else
"110111011111" when X = 258 AND Y = 29 else
"110111011111" when X = 259 AND Y = 29 else
"110111011111" when X = 260 AND Y = 29 else
"110111011111" when X = 261 AND Y = 29 else
"110111011111" when X = 262 AND Y = 29 else
"110111011111" when X = 263 AND Y = 29 else
"110111011111" when X = 264 AND Y = 29 else
"110111011111" when X = 265 AND Y = 29 else
"110111011111" when X = 266 AND Y = 29 else
"110111011111" when X = 267 AND Y = 29 else
"110111011111" when X = 268 AND Y = 29 else
"110111011111" when X = 269 AND Y = 29 else
"110111011111" when X = 270 AND Y = 29 else
"110111011111" when X = 271 AND Y = 29 else
"110111011111" when X = 272 AND Y = 29 else
"110111011111" when X = 273 AND Y = 29 else
"110111011111" when X = 274 AND Y = 29 else
"110111011111" when X = 275 AND Y = 29 else
"110111011111" when X = 276 AND Y = 29 else
"110111011111" when X = 277 AND Y = 29 else
"110111011111" when X = 278 AND Y = 29 else
"110111011111" when X = 279 AND Y = 29 else
"000000000000" when X = 280 AND Y = 29 else
"000000000000" when X = 281 AND Y = 29 else
"000000000000" when X = 282 AND Y = 29 else
"000000000000" when X = 283 AND Y = 29 else
"000000000000" when X = 284 AND Y = 29 else
"000000000000" when X = 285 AND Y = 29 else
"000000000000" when X = 286 AND Y = 29 else
"000000000000" when X = 287 AND Y = 29 else
"000000000000" when X = 288 AND Y = 29 else
"000000000000" when X = 289 AND Y = 29 else
"000000000000" when X = 290 AND Y = 29 else
"000000000000" when X = 291 AND Y = 29 else
"000000000000" when X = 292 AND Y = 29 else
"000000000000" when X = 293 AND Y = 29 else
"000000000000" when X = 294 AND Y = 29 else
"000000000000" when X = 295 AND Y = 29 else
"000000000000" when X = 296 AND Y = 29 else
"000000000000" when X = 297 AND Y = 29 else
"000000000000" when X = 298 AND Y = 29 else
"000000000000" when X = 299 AND Y = 29 else
"000000000000" when X = 300 AND Y = 29 else
"000000000000" when X = 301 AND Y = 29 else
"000000000000" when X = 302 AND Y = 29 else
"000000000000" when X = 303 AND Y = 29 else
"000000000000" when X = 304 AND Y = 29 else
"000000000000" when X = 305 AND Y = 29 else
"000000000000" when X = 306 AND Y = 29 else
"000000000000" when X = 307 AND Y = 29 else
"000000000000" when X = 308 AND Y = 29 else
"000000000000" when X = 309 AND Y = 29 else
"000000000000" when X = 310 AND Y = 29 else
"000000000000" when X = 311 AND Y = 29 else
"000000000000" when X = 312 AND Y = 29 else
"000000000000" when X = 313 AND Y = 29 else
"000000000000" when X = 314 AND Y = 29 else
"000000000000" when X = 315 AND Y = 29 else
"000000000000" when X = 316 AND Y = 29 else
"000000000000" when X = 317 AND Y = 29 else
"000000000000" when X = 318 AND Y = 29 else
"000000000000" when X = 319 AND Y = 29 else
"000000000000" when X = 320 AND Y = 29 else
"000000000000" when X = 321 AND Y = 29 else
"000000000000" when X = 322 AND Y = 29 else
"000000000000" when X = 323 AND Y = 29 else
"000000000000" when X = 324 AND Y = 29 else
"000000000000" when X = 0 AND Y = 30 else
"000000000000" when X = 1 AND Y = 30 else
"000000000000" when X = 2 AND Y = 30 else
"000000000000" when X = 3 AND Y = 30 else
"000000000000" when X = 4 AND Y = 30 else
"000000000000" when X = 5 AND Y = 30 else
"000000000000" when X = 6 AND Y = 30 else
"000000000000" when X = 7 AND Y = 30 else
"000000000000" when X = 8 AND Y = 30 else
"000000000000" when X = 9 AND Y = 30 else
"000000000000" when X = 10 AND Y = 30 else
"000000000000" when X = 11 AND Y = 30 else
"000000000000" when X = 12 AND Y = 30 else
"000000000000" when X = 13 AND Y = 30 else
"000000000000" when X = 14 AND Y = 30 else
"000000000000" when X = 15 AND Y = 30 else
"000000000000" when X = 16 AND Y = 30 else
"000000000000" when X = 17 AND Y = 30 else
"000000000000" when X = 18 AND Y = 30 else
"000000000000" when X = 19 AND Y = 30 else
"000000000000" when X = 20 AND Y = 30 else
"000000000000" when X = 21 AND Y = 30 else
"000000000000" when X = 22 AND Y = 30 else
"000000000000" when X = 23 AND Y = 30 else
"000000000000" when X = 24 AND Y = 30 else
"000000000000" when X = 25 AND Y = 30 else
"000000000000" when X = 26 AND Y = 30 else
"000000000000" when X = 27 AND Y = 30 else
"000000000000" when X = 28 AND Y = 30 else
"000000000000" when X = 29 AND Y = 30 else
"000000000000" when X = 30 AND Y = 30 else
"000000000000" when X = 31 AND Y = 30 else
"000000000000" when X = 32 AND Y = 30 else
"000000000000" when X = 33 AND Y = 30 else
"000000000000" when X = 34 AND Y = 30 else
"000000000000" when X = 35 AND Y = 30 else
"000000000000" when X = 36 AND Y = 30 else
"000000000000" when X = 37 AND Y = 30 else
"000000000000" when X = 38 AND Y = 30 else
"000000000000" when X = 39 AND Y = 30 else
"100010011101" when X = 40 AND Y = 30 else
"100010011101" when X = 41 AND Y = 30 else
"100010011101" when X = 42 AND Y = 30 else
"100010011101" when X = 43 AND Y = 30 else
"100010011101" when X = 44 AND Y = 30 else
"100010011101" when X = 45 AND Y = 30 else
"100010011101" when X = 46 AND Y = 30 else
"100010011101" when X = 47 AND Y = 30 else
"100010011101" when X = 48 AND Y = 30 else
"100010011101" when X = 49 AND Y = 30 else
"110111011111" when X = 50 AND Y = 30 else
"110111011111" when X = 51 AND Y = 30 else
"110111011111" when X = 52 AND Y = 30 else
"110111011111" when X = 53 AND Y = 30 else
"110111011111" when X = 54 AND Y = 30 else
"110111011111" when X = 55 AND Y = 30 else
"110111011111" when X = 56 AND Y = 30 else
"110111011111" when X = 57 AND Y = 30 else
"110111011111" when X = 58 AND Y = 30 else
"110111011111" when X = 59 AND Y = 30 else
"111111111111" when X = 60 AND Y = 30 else
"111111111111" when X = 61 AND Y = 30 else
"111111111111" when X = 62 AND Y = 30 else
"111111111111" when X = 63 AND Y = 30 else
"111111111111" when X = 64 AND Y = 30 else
"111111111111" when X = 65 AND Y = 30 else
"111111111111" when X = 66 AND Y = 30 else
"111111111111" when X = 67 AND Y = 30 else
"111111111111" when X = 68 AND Y = 30 else
"111111111111" when X = 69 AND Y = 30 else
"111111111111" when X = 70 AND Y = 30 else
"111111111111" when X = 71 AND Y = 30 else
"111111111111" when X = 72 AND Y = 30 else
"111111111111" when X = 73 AND Y = 30 else
"111111111111" when X = 74 AND Y = 30 else
"111111111111" when X = 75 AND Y = 30 else
"111111111111" when X = 76 AND Y = 30 else
"111111111111" when X = 77 AND Y = 30 else
"111111111111" when X = 78 AND Y = 30 else
"111111111111" when X = 79 AND Y = 30 else
"111111111111" when X = 80 AND Y = 30 else
"111111111111" when X = 81 AND Y = 30 else
"111111111111" when X = 82 AND Y = 30 else
"111111111111" when X = 83 AND Y = 30 else
"111111111111" when X = 84 AND Y = 30 else
"111111111111" when X = 85 AND Y = 30 else
"111111111111" when X = 86 AND Y = 30 else
"111111111111" when X = 87 AND Y = 30 else
"111111111111" when X = 88 AND Y = 30 else
"111111111111" when X = 89 AND Y = 30 else
"111111111111" when X = 90 AND Y = 30 else
"111111111111" when X = 91 AND Y = 30 else
"111111111111" when X = 92 AND Y = 30 else
"111111111111" when X = 93 AND Y = 30 else
"111111111111" when X = 94 AND Y = 30 else
"111111111111" when X = 95 AND Y = 30 else
"111111111111" when X = 96 AND Y = 30 else
"111111111111" when X = 97 AND Y = 30 else
"111111111111" when X = 98 AND Y = 30 else
"111111111111" when X = 99 AND Y = 30 else
"111111111111" when X = 100 AND Y = 30 else
"111111111111" when X = 101 AND Y = 30 else
"111111111111" when X = 102 AND Y = 30 else
"111111111111" when X = 103 AND Y = 30 else
"111111111111" when X = 104 AND Y = 30 else
"111111111111" when X = 105 AND Y = 30 else
"111111111111" when X = 106 AND Y = 30 else
"111111111111" when X = 107 AND Y = 30 else
"111111111111" when X = 108 AND Y = 30 else
"111111111111" when X = 109 AND Y = 30 else
"111111111111" when X = 110 AND Y = 30 else
"111111111111" when X = 111 AND Y = 30 else
"111111111111" when X = 112 AND Y = 30 else
"111111111111" when X = 113 AND Y = 30 else
"111111111111" when X = 114 AND Y = 30 else
"111111111111" when X = 115 AND Y = 30 else
"111111111111" when X = 116 AND Y = 30 else
"111111111111" when X = 117 AND Y = 30 else
"111111111111" when X = 118 AND Y = 30 else
"111111111111" when X = 119 AND Y = 30 else
"111111111111" when X = 120 AND Y = 30 else
"111111111111" when X = 121 AND Y = 30 else
"111111111111" when X = 122 AND Y = 30 else
"111111111111" when X = 123 AND Y = 30 else
"111111111111" when X = 124 AND Y = 30 else
"111111111111" when X = 125 AND Y = 30 else
"111111111111" when X = 126 AND Y = 30 else
"111111111111" when X = 127 AND Y = 30 else
"111111111111" when X = 128 AND Y = 30 else
"111111111111" when X = 129 AND Y = 30 else
"111111111111" when X = 130 AND Y = 30 else
"111111111111" when X = 131 AND Y = 30 else
"111111111111" when X = 132 AND Y = 30 else
"111111111111" when X = 133 AND Y = 30 else
"111111111111" when X = 134 AND Y = 30 else
"111111111111" when X = 135 AND Y = 30 else
"111111111111" when X = 136 AND Y = 30 else
"111111111111" when X = 137 AND Y = 30 else
"111111111111" when X = 138 AND Y = 30 else
"111111111111" when X = 139 AND Y = 30 else
"111111111111" when X = 140 AND Y = 30 else
"111111111111" when X = 141 AND Y = 30 else
"111111111111" when X = 142 AND Y = 30 else
"111111111111" when X = 143 AND Y = 30 else
"111111111111" when X = 144 AND Y = 30 else
"111111111111" when X = 145 AND Y = 30 else
"111111111111" when X = 146 AND Y = 30 else
"111111111111" when X = 147 AND Y = 30 else
"111111111111" when X = 148 AND Y = 30 else
"111111111111" when X = 149 AND Y = 30 else
"111111111111" when X = 150 AND Y = 30 else
"111111111111" when X = 151 AND Y = 30 else
"111111111111" when X = 152 AND Y = 30 else
"111111111111" when X = 153 AND Y = 30 else
"111111111111" when X = 154 AND Y = 30 else
"111111111111" when X = 155 AND Y = 30 else
"111111111111" when X = 156 AND Y = 30 else
"111111111111" when X = 157 AND Y = 30 else
"111111111111" when X = 158 AND Y = 30 else
"111111111111" when X = 159 AND Y = 30 else
"111111111111" when X = 160 AND Y = 30 else
"111111111111" when X = 161 AND Y = 30 else
"111111111111" when X = 162 AND Y = 30 else
"111111111111" when X = 163 AND Y = 30 else
"111111111111" when X = 164 AND Y = 30 else
"111111111111" when X = 165 AND Y = 30 else
"111111111111" when X = 166 AND Y = 30 else
"111111111111" when X = 167 AND Y = 30 else
"111111111111" when X = 168 AND Y = 30 else
"111111111111" when X = 169 AND Y = 30 else
"111111111111" when X = 170 AND Y = 30 else
"111111111111" when X = 171 AND Y = 30 else
"111111111111" when X = 172 AND Y = 30 else
"111111111111" when X = 173 AND Y = 30 else
"111111111111" when X = 174 AND Y = 30 else
"111111111111" when X = 175 AND Y = 30 else
"111111111111" when X = 176 AND Y = 30 else
"111111111111" when X = 177 AND Y = 30 else
"111111111111" when X = 178 AND Y = 30 else
"111111111111" when X = 179 AND Y = 30 else
"111111111111" when X = 180 AND Y = 30 else
"111111111111" when X = 181 AND Y = 30 else
"111111111111" when X = 182 AND Y = 30 else
"111111111111" when X = 183 AND Y = 30 else
"111111111111" when X = 184 AND Y = 30 else
"111111111111" when X = 185 AND Y = 30 else
"111111111111" when X = 186 AND Y = 30 else
"111111111111" when X = 187 AND Y = 30 else
"111111111111" when X = 188 AND Y = 30 else
"111111111111" when X = 189 AND Y = 30 else
"000000000000" when X = 190 AND Y = 30 else
"000000000000" when X = 191 AND Y = 30 else
"000000000000" when X = 192 AND Y = 30 else
"000000000000" when X = 193 AND Y = 30 else
"000000000000" when X = 194 AND Y = 30 else
"000000000000" when X = 195 AND Y = 30 else
"000000000000" when X = 196 AND Y = 30 else
"000000000000" when X = 197 AND Y = 30 else
"000000000000" when X = 198 AND Y = 30 else
"000000000000" when X = 199 AND Y = 30 else
"000000000000" when X = 200 AND Y = 30 else
"000000000000" when X = 201 AND Y = 30 else
"000000000000" when X = 202 AND Y = 30 else
"000000000000" when X = 203 AND Y = 30 else
"000000000000" when X = 204 AND Y = 30 else
"000000000000" when X = 205 AND Y = 30 else
"000000000000" when X = 206 AND Y = 30 else
"000000000000" when X = 207 AND Y = 30 else
"000000000000" when X = 208 AND Y = 30 else
"000000000000" when X = 209 AND Y = 30 else
"000000000000" when X = 210 AND Y = 30 else
"000000000000" when X = 211 AND Y = 30 else
"000000000000" when X = 212 AND Y = 30 else
"000000000000" when X = 213 AND Y = 30 else
"000000000000" when X = 214 AND Y = 30 else
"000000000000" when X = 215 AND Y = 30 else
"000000000000" when X = 216 AND Y = 30 else
"000000000000" when X = 217 AND Y = 30 else
"000000000000" when X = 218 AND Y = 30 else
"000000000000" when X = 219 AND Y = 30 else
"000000000000" when X = 220 AND Y = 30 else
"000000000000" when X = 221 AND Y = 30 else
"000000000000" when X = 222 AND Y = 30 else
"000000000000" when X = 223 AND Y = 30 else
"000000000000" when X = 224 AND Y = 30 else
"111111111111" when X = 225 AND Y = 30 else
"111111111111" when X = 226 AND Y = 30 else
"111111111111" when X = 227 AND Y = 30 else
"111111111111" when X = 228 AND Y = 30 else
"111111111111" when X = 229 AND Y = 30 else
"111111111111" when X = 230 AND Y = 30 else
"111111111111" when X = 231 AND Y = 30 else
"111111111111" when X = 232 AND Y = 30 else
"111111111111" when X = 233 AND Y = 30 else
"111111111111" when X = 234 AND Y = 30 else
"111111111111" when X = 235 AND Y = 30 else
"111111111111" when X = 236 AND Y = 30 else
"111111111111" when X = 237 AND Y = 30 else
"111111111111" when X = 238 AND Y = 30 else
"111111111111" when X = 239 AND Y = 30 else
"111111111111" when X = 240 AND Y = 30 else
"111111111111" when X = 241 AND Y = 30 else
"111111111111" when X = 242 AND Y = 30 else
"111111111111" when X = 243 AND Y = 30 else
"111111111111" when X = 244 AND Y = 30 else
"111111111111" when X = 245 AND Y = 30 else
"111111111111" when X = 246 AND Y = 30 else
"111111111111" when X = 247 AND Y = 30 else
"111111111111" when X = 248 AND Y = 30 else
"111111111111" when X = 249 AND Y = 30 else
"111111111111" when X = 250 AND Y = 30 else
"111111111111" when X = 251 AND Y = 30 else
"111111111111" when X = 252 AND Y = 30 else
"111111111111" when X = 253 AND Y = 30 else
"111111111111" when X = 254 AND Y = 30 else
"110111011111" when X = 255 AND Y = 30 else
"110111011111" when X = 256 AND Y = 30 else
"110111011111" when X = 257 AND Y = 30 else
"110111011111" when X = 258 AND Y = 30 else
"110111011111" when X = 259 AND Y = 30 else
"110111011111" when X = 260 AND Y = 30 else
"110111011111" when X = 261 AND Y = 30 else
"110111011111" when X = 262 AND Y = 30 else
"110111011111" when X = 263 AND Y = 30 else
"110111011111" when X = 264 AND Y = 30 else
"110111011111" when X = 265 AND Y = 30 else
"110111011111" when X = 266 AND Y = 30 else
"110111011111" when X = 267 AND Y = 30 else
"110111011111" when X = 268 AND Y = 30 else
"110111011111" when X = 269 AND Y = 30 else
"110111011111" when X = 270 AND Y = 30 else
"110111011111" when X = 271 AND Y = 30 else
"110111011111" when X = 272 AND Y = 30 else
"110111011111" when X = 273 AND Y = 30 else
"110111011111" when X = 274 AND Y = 30 else
"110111011111" when X = 275 AND Y = 30 else
"110111011111" when X = 276 AND Y = 30 else
"110111011111" when X = 277 AND Y = 30 else
"110111011111" when X = 278 AND Y = 30 else
"110111011111" when X = 279 AND Y = 30 else
"000000000000" when X = 280 AND Y = 30 else
"000000000000" when X = 281 AND Y = 30 else
"000000000000" when X = 282 AND Y = 30 else
"000000000000" when X = 283 AND Y = 30 else
"000000000000" when X = 284 AND Y = 30 else
"000000000000" when X = 285 AND Y = 30 else
"000000000000" when X = 286 AND Y = 30 else
"000000000000" when X = 287 AND Y = 30 else
"000000000000" when X = 288 AND Y = 30 else
"000000000000" when X = 289 AND Y = 30 else
"000000000000" when X = 290 AND Y = 30 else
"000000000000" when X = 291 AND Y = 30 else
"000000000000" when X = 292 AND Y = 30 else
"000000000000" when X = 293 AND Y = 30 else
"000000000000" when X = 294 AND Y = 30 else
"000000000000" when X = 295 AND Y = 30 else
"000000000000" when X = 296 AND Y = 30 else
"000000000000" when X = 297 AND Y = 30 else
"000000000000" when X = 298 AND Y = 30 else
"000000000000" when X = 299 AND Y = 30 else
"000000000000" when X = 300 AND Y = 30 else
"000000000000" when X = 301 AND Y = 30 else
"000000000000" when X = 302 AND Y = 30 else
"000000000000" when X = 303 AND Y = 30 else
"000000000000" when X = 304 AND Y = 30 else
"000000000000" when X = 305 AND Y = 30 else
"000000000000" when X = 306 AND Y = 30 else
"000000000000" when X = 307 AND Y = 30 else
"000000000000" when X = 308 AND Y = 30 else
"000000000000" when X = 309 AND Y = 30 else
"000000000000" when X = 310 AND Y = 30 else
"000000000000" when X = 311 AND Y = 30 else
"000000000000" when X = 312 AND Y = 30 else
"000000000000" when X = 313 AND Y = 30 else
"000000000000" when X = 314 AND Y = 30 else
"000000000000" when X = 315 AND Y = 30 else
"000000000000" when X = 316 AND Y = 30 else
"000000000000" when X = 317 AND Y = 30 else
"000000000000" when X = 318 AND Y = 30 else
"000000000000" when X = 319 AND Y = 30 else
"000000000000" when X = 320 AND Y = 30 else
"000000000000" when X = 321 AND Y = 30 else
"000000000000" when X = 322 AND Y = 30 else
"000000000000" when X = 323 AND Y = 30 else
"000000000000" when X = 324 AND Y = 30 else
"000000000000" when X = 0 AND Y = 31 else
"000000000000" when X = 1 AND Y = 31 else
"000000000000" when X = 2 AND Y = 31 else
"000000000000" when X = 3 AND Y = 31 else
"000000000000" when X = 4 AND Y = 31 else
"000000000000" when X = 5 AND Y = 31 else
"000000000000" when X = 6 AND Y = 31 else
"000000000000" when X = 7 AND Y = 31 else
"000000000000" when X = 8 AND Y = 31 else
"000000000000" when X = 9 AND Y = 31 else
"000000000000" when X = 10 AND Y = 31 else
"000000000000" when X = 11 AND Y = 31 else
"000000000000" when X = 12 AND Y = 31 else
"000000000000" when X = 13 AND Y = 31 else
"000000000000" when X = 14 AND Y = 31 else
"000000000000" when X = 15 AND Y = 31 else
"000000000000" when X = 16 AND Y = 31 else
"000000000000" when X = 17 AND Y = 31 else
"000000000000" when X = 18 AND Y = 31 else
"000000000000" when X = 19 AND Y = 31 else
"000000000000" when X = 20 AND Y = 31 else
"000000000000" when X = 21 AND Y = 31 else
"000000000000" when X = 22 AND Y = 31 else
"000000000000" when X = 23 AND Y = 31 else
"000000000000" when X = 24 AND Y = 31 else
"000000000000" when X = 25 AND Y = 31 else
"000000000000" when X = 26 AND Y = 31 else
"000000000000" when X = 27 AND Y = 31 else
"000000000000" when X = 28 AND Y = 31 else
"000000000000" when X = 29 AND Y = 31 else
"000000000000" when X = 30 AND Y = 31 else
"000000000000" when X = 31 AND Y = 31 else
"000000000000" when X = 32 AND Y = 31 else
"000000000000" when X = 33 AND Y = 31 else
"000000000000" when X = 34 AND Y = 31 else
"000000000000" when X = 35 AND Y = 31 else
"000000000000" when X = 36 AND Y = 31 else
"000000000000" when X = 37 AND Y = 31 else
"000000000000" when X = 38 AND Y = 31 else
"000000000000" when X = 39 AND Y = 31 else
"100010011101" when X = 40 AND Y = 31 else
"100010011101" when X = 41 AND Y = 31 else
"100010011101" when X = 42 AND Y = 31 else
"100010011101" when X = 43 AND Y = 31 else
"100010011101" when X = 44 AND Y = 31 else
"100010011101" when X = 45 AND Y = 31 else
"100010011101" when X = 46 AND Y = 31 else
"100010011101" when X = 47 AND Y = 31 else
"100010011101" when X = 48 AND Y = 31 else
"100010011101" when X = 49 AND Y = 31 else
"110111011111" when X = 50 AND Y = 31 else
"110111011111" when X = 51 AND Y = 31 else
"110111011111" when X = 52 AND Y = 31 else
"110111011111" when X = 53 AND Y = 31 else
"110111011111" when X = 54 AND Y = 31 else
"110111011111" when X = 55 AND Y = 31 else
"110111011111" when X = 56 AND Y = 31 else
"110111011111" when X = 57 AND Y = 31 else
"110111011111" when X = 58 AND Y = 31 else
"110111011111" when X = 59 AND Y = 31 else
"111111111111" when X = 60 AND Y = 31 else
"111111111111" when X = 61 AND Y = 31 else
"111111111111" when X = 62 AND Y = 31 else
"111111111111" when X = 63 AND Y = 31 else
"111111111111" when X = 64 AND Y = 31 else
"111111111111" when X = 65 AND Y = 31 else
"111111111111" when X = 66 AND Y = 31 else
"111111111111" when X = 67 AND Y = 31 else
"111111111111" when X = 68 AND Y = 31 else
"111111111111" when X = 69 AND Y = 31 else
"111111111111" when X = 70 AND Y = 31 else
"111111111111" when X = 71 AND Y = 31 else
"111111111111" when X = 72 AND Y = 31 else
"111111111111" when X = 73 AND Y = 31 else
"111111111111" when X = 74 AND Y = 31 else
"111111111111" when X = 75 AND Y = 31 else
"111111111111" when X = 76 AND Y = 31 else
"111111111111" when X = 77 AND Y = 31 else
"111111111111" when X = 78 AND Y = 31 else
"111111111111" when X = 79 AND Y = 31 else
"111111111111" when X = 80 AND Y = 31 else
"111111111111" when X = 81 AND Y = 31 else
"111111111111" when X = 82 AND Y = 31 else
"111111111111" when X = 83 AND Y = 31 else
"111111111111" when X = 84 AND Y = 31 else
"111111111111" when X = 85 AND Y = 31 else
"111111111111" when X = 86 AND Y = 31 else
"111111111111" when X = 87 AND Y = 31 else
"111111111111" when X = 88 AND Y = 31 else
"111111111111" when X = 89 AND Y = 31 else
"111111111111" when X = 90 AND Y = 31 else
"111111111111" when X = 91 AND Y = 31 else
"111111111111" when X = 92 AND Y = 31 else
"111111111111" when X = 93 AND Y = 31 else
"111111111111" when X = 94 AND Y = 31 else
"111111111111" when X = 95 AND Y = 31 else
"111111111111" when X = 96 AND Y = 31 else
"111111111111" when X = 97 AND Y = 31 else
"111111111111" when X = 98 AND Y = 31 else
"111111111111" when X = 99 AND Y = 31 else
"111111111111" when X = 100 AND Y = 31 else
"111111111111" when X = 101 AND Y = 31 else
"111111111111" when X = 102 AND Y = 31 else
"111111111111" when X = 103 AND Y = 31 else
"111111111111" when X = 104 AND Y = 31 else
"111111111111" when X = 105 AND Y = 31 else
"111111111111" when X = 106 AND Y = 31 else
"111111111111" when X = 107 AND Y = 31 else
"111111111111" when X = 108 AND Y = 31 else
"111111111111" when X = 109 AND Y = 31 else
"111111111111" when X = 110 AND Y = 31 else
"111111111111" when X = 111 AND Y = 31 else
"111111111111" when X = 112 AND Y = 31 else
"111111111111" when X = 113 AND Y = 31 else
"111111111111" when X = 114 AND Y = 31 else
"111111111111" when X = 115 AND Y = 31 else
"111111111111" when X = 116 AND Y = 31 else
"111111111111" when X = 117 AND Y = 31 else
"111111111111" when X = 118 AND Y = 31 else
"111111111111" when X = 119 AND Y = 31 else
"111111111111" when X = 120 AND Y = 31 else
"111111111111" when X = 121 AND Y = 31 else
"111111111111" when X = 122 AND Y = 31 else
"111111111111" when X = 123 AND Y = 31 else
"111111111111" when X = 124 AND Y = 31 else
"111111111111" when X = 125 AND Y = 31 else
"111111111111" when X = 126 AND Y = 31 else
"111111111111" when X = 127 AND Y = 31 else
"111111111111" when X = 128 AND Y = 31 else
"111111111111" when X = 129 AND Y = 31 else
"111111111111" when X = 130 AND Y = 31 else
"111111111111" when X = 131 AND Y = 31 else
"111111111111" when X = 132 AND Y = 31 else
"111111111111" when X = 133 AND Y = 31 else
"111111111111" when X = 134 AND Y = 31 else
"111111111111" when X = 135 AND Y = 31 else
"111111111111" when X = 136 AND Y = 31 else
"111111111111" when X = 137 AND Y = 31 else
"111111111111" when X = 138 AND Y = 31 else
"111111111111" when X = 139 AND Y = 31 else
"111111111111" when X = 140 AND Y = 31 else
"111111111111" when X = 141 AND Y = 31 else
"111111111111" when X = 142 AND Y = 31 else
"111111111111" when X = 143 AND Y = 31 else
"111111111111" when X = 144 AND Y = 31 else
"111111111111" when X = 145 AND Y = 31 else
"111111111111" when X = 146 AND Y = 31 else
"111111111111" when X = 147 AND Y = 31 else
"111111111111" when X = 148 AND Y = 31 else
"111111111111" when X = 149 AND Y = 31 else
"111111111111" when X = 150 AND Y = 31 else
"111111111111" when X = 151 AND Y = 31 else
"111111111111" when X = 152 AND Y = 31 else
"111111111111" when X = 153 AND Y = 31 else
"111111111111" when X = 154 AND Y = 31 else
"111111111111" when X = 155 AND Y = 31 else
"111111111111" when X = 156 AND Y = 31 else
"111111111111" when X = 157 AND Y = 31 else
"111111111111" when X = 158 AND Y = 31 else
"111111111111" when X = 159 AND Y = 31 else
"111111111111" when X = 160 AND Y = 31 else
"111111111111" when X = 161 AND Y = 31 else
"111111111111" when X = 162 AND Y = 31 else
"111111111111" when X = 163 AND Y = 31 else
"111111111111" when X = 164 AND Y = 31 else
"111111111111" when X = 165 AND Y = 31 else
"111111111111" when X = 166 AND Y = 31 else
"111111111111" when X = 167 AND Y = 31 else
"111111111111" when X = 168 AND Y = 31 else
"111111111111" when X = 169 AND Y = 31 else
"111111111111" when X = 170 AND Y = 31 else
"111111111111" when X = 171 AND Y = 31 else
"111111111111" when X = 172 AND Y = 31 else
"111111111111" when X = 173 AND Y = 31 else
"111111111111" when X = 174 AND Y = 31 else
"111111111111" when X = 175 AND Y = 31 else
"111111111111" when X = 176 AND Y = 31 else
"111111111111" when X = 177 AND Y = 31 else
"111111111111" when X = 178 AND Y = 31 else
"111111111111" when X = 179 AND Y = 31 else
"111111111111" when X = 180 AND Y = 31 else
"111111111111" when X = 181 AND Y = 31 else
"111111111111" when X = 182 AND Y = 31 else
"111111111111" when X = 183 AND Y = 31 else
"111111111111" when X = 184 AND Y = 31 else
"111111111111" when X = 185 AND Y = 31 else
"111111111111" when X = 186 AND Y = 31 else
"111111111111" when X = 187 AND Y = 31 else
"111111111111" when X = 188 AND Y = 31 else
"111111111111" when X = 189 AND Y = 31 else
"000000000000" when X = 190 AND Y = 31 else
"000000000000" when X = 191 AND Y = 31 else
"000000000000" when X = 192 AND Y = 31 else
"000000000000" when X = 193 AND Y = 31 else
"000000000000" when X = 194 AND Y = 31 else
"000000000000" when X = 195 AND Y = 31 else
"000000000000" when X = 196 AND Y = 31 else
"000000000000" when X = 197 AND Y = 31 else
"000000000000" when X = 198 AND Y = 31 else
"000000000000" when X = 199 AND Y = 31 else
"000000000000" when X = 200 AND Y = 31 else
"000000000000" when X = 201 AND Y = 31 else
"000000000000" when X = 202 AND Y = 31 else
"000000000000" when X = 203 AND Y = 31 else
"000000000000" when X = 204 AND Y = 31 else
"000000000000" when X = 205 AND Y = 31 else
"000000000000" when X = 206 AND Y = 31 else
"000000000000" when X = 207 AND Y = 31 else
"000000000000" when X = 208 AND Y = 31 else
"000000000000" when X = 209 AND Y = 31 else
"000000000000" when X = 210 AND Y = 31 else
"000000000000" when X = 211 AND Y = 31 else
"000000000000" when X = 212 AND Y = 31 else
"000000000000" when X = 213 AND Y = 31 else
"000000000000" when X = 214 AND Y = 31 else
"000000000000" when X = 215 AND Y = 31 else
"000000000000" when X = 216 AND Y = 31 else
"000000000000" when X = 217 AND Y = 31 else
"000000000000" when X = 218 AND Y = 31 else
"000000000000" when X = 219 AND Y = 31 else
"000000000000" when X = 220 AND Y = 31 else
"000000000000" when X = 221 AND Y = 31 else
"000000000000" when X = 222 AND Y = 31 else
"000000000000" when X = 223 AND Y = 31 else
"000000000000" when X = 224 AND Y = 31 else
"111111111111" when X = 225 AND Y = 31 else
"111111111111" when X = 226 AND Y = 31 else
"111111111111" when X = 227 AND Y = 31 else
"111111111111" when X = 228 AND Y = 31 else
"111111111111" when X = 229 AND Y = 31 else
"111111111111" when X = 230 AND Y = 31 else
"111111111111" when X = 231 AND Y = 31 else
"111111111111" when X = 232 AND Y = 31 else
"111111111111" when X = 233 AND Y = 31 else
"111111111111" when X = 234 AND Y = 31 else
"111111111111" when X = 235 AND Y = 31 else
"111111111111" when X = 236 AND Y = 31 else
"111111111111" when X = 237 AND Y = 31 else
"111111111111" when X = 238 AND Y = 31 else
"111111111111" when X = 239 AND Y = 31 else
"111111111111" when X = 240 AND Y = 31 else
"111111111111" when X = 241 AND Y = 31 else
"111111111111" when X = 242 AND Y = 31 else
"111111111111" when X = 243 AND Y = 31 else
"111111111111" when X = 244 AND Y = 31 else
"111111111111" when X = 245 AND Y = 31 else
"111111111111" when X = 246 AND Y = 31 else
"111111111111" when X = 247 AND Y = 31 else
"111111111111" when X = 248 AND Y = 31 else
"111111111111" when X = 249 AND Y = 31 else
"111111111111" when X = 250 AND Y = 31 else
"111111111111" when X = 251 AND Y = 31 else
"111111111111" when X = 252 AND Y = 31 else
"111111111111" when X = 253 AND Y = 31 else
"111111111111" when X = 254 AND Y = 31 else
"110111011111" when X = 255 AND Y = 31 else
"110111011111" when X = 256 AND Y = 31 else
"110111011111" when X = 257 AND Y = 31 else
"110111011111" when X = 258 AND Y = 31 else
"110111011111" when X = 259 AND Y = 31 else
"110111011111" when X = 260 AND Y = 31 else
"110111011111" when X = 261 AND Y = 31 else
"110111011111" when X = 262 AND Y = 31 else
"110111011111" when X = 263 AND Y = 31 else
"110111011111" when X = 264 AND Y = 31 else
"110111011111" when X = 265 AND Y = 31 else
"110111011111" when X = 266 AND Y = 31 else
"110111011111" when X = 267 AND Y = 31 else
"110111011111" when X = 268 AND Y = 31 else
"110111011111" when X = 269 AND Y = 31 else
"110111011111" when X = 270 AND Y = 31 else
"110111011111" when X = 271 AND Y = 31 else
"110111011111" when X = 272 AND Y = 31 else
"110111011111" when X = 273 AND Y = 31 else
"110111011111" when X = 274 AND Y = 31 else
"110111011111" when X = 275 AND Y = 31 else
"110111011111" when X = 276 AND Y = 31 else
"110111011111" when X = 277 AND Y = 31 else
"110111011111" when X = 278 AND Y = 31 else
"110111011111" when X = 279 AND Y = 31 else
"000000000000" when X = 280 AND Y = 31 else
"000000000000" when X = 281 AND Y = 31 else
"000000000000" when X = 282 AND Y = 31 else
"000000000000" when X = 283 AND Y = 31 else
"000000000000" when X = 284 AND Y = 31 else
"000000000000" when X = 285 AND Y = 31 else
"000000000000" when X = 286 AND Y = 31 else
"000000000000" when X = 287 AND Y = 31 else
"000000000000" when X = 288 AND Y = 31 else
"000000000000" when X = 289 AND Y = 31 else
"000000000000" when X = 290 AND Y = 31 else
"000000000000" when X = 291 AND Y = 31 else
"000000000000" when X = 292 AND Y = 31 else
"000000000000" when X = 293 AND Y = 31 else
"000000000000" when X = 294 AND Y = 31 else
"000000000000" when X = 295 AND Y = 31 else
"000000000000" when X = 296 AND Y = 31 else
"000000000000" when X = 297 AND Y = 31 else
"000000000000" when X = 298 AND Y = 31 else
"000000000000" when X = 299 AND Y = 31 else
"000000000000" when X = 300 AND Y = 31 else
"000000000000" when X = 301 AND Y = 31 else
"000000000000" when X = 302 AND Y = 31 else
"000000000000" when X = 303 AND Y = 31 else
"000000000000" when X = 304 AND Y = 31 else
"000000000000" when X = 305 AND Y = 31 else
"000000000000" when X = 306 AND Y = 31 else
"000000000000" when X = 307 AND Y = 31 else
"000000000000" when X = 308 AND Y = 31 else
"000000000000" when X = 309 AND Y = 31 else
"000000000000" when X = 310 AND Y = 31 else
"000000000000" when X = 311 AND Y = 31 else
"000000000000" when X = 312 AND Y = 31 else
"000000000000" when X = 313 AND Y = 31 else
"000000000000" when X = 314 AND Y = 31 else
"000000000000" when X = 315 AND Y = 31 else
"000000000000" when X = 316 AND Y = 31 else
"000000000000" when X = 317 AND Y = 31 else
"000000000000" when X = 318 AND Y = 31 else
"000000000000" when X = 319 AND Y = 31 else
"000000000000" when X = 320 AND Y = 31 else
"000000000000" when X = 321 AND Y = 31 else
"000000000000" when X = 322 AND Y = 31 else
"000000000000" when X = 323 AND Y = 31 else
"000000000000" when X = 324 AND Y = 31 else
"000000000000" when X = 0 AND Y = 32 else
"000000000000" when X = 1 AND Y = 32 else
"000000000000" when X = 2 AND Y = 32 else
"000000000000" when X = 3 AND Y = 32 else
"000000000000" when X = 4 AND Y = 32 else
"000000000000" when X = 5 AND Y = 32 else
"000000000000" when X = 6 AND Y = 32 else
"000000000000" when X = 7 AND Y = 32 else
"000000000000" when X = 8 AND Y = 32 else
"000000000000" when X = 9 AND Y = 32 else
"000000000000" when X = 10 AND Y = 32 else
"000000000000" when X = 11 AND Y = 32 else
"000000000000" when X = 12 AND Y = 32 else
"000000000000" when X = 13 AND Y = 32 else
"000000000000" when X = 14 AND Y = 32 else
"000000000000" when X = 15 AND Y = 32 else
"000000000000" when X = 16 AND Y = 32 else
"000000000000" when X = 17 AND Y = 32 else
"000000000000" when X = 18 AND Y = 32 else
"000000000000" when X = 19 AND Y = 32 else
"000000000000" when X = 20 AND Y = 32 else
"000000000000" when X = 21 AND Y = 32 else
"000000000000" when X = 22 AND Y = 32 else
"000000000000" when X = 23 AND Y = 32 else
"000000000000" when X = 24 AND Y = 32 else
"000000000000" when X = 25 AND Y = 32 else
"000000000000" when X = 26 AND Y = 32 else
"000000000000" when X = 27 AND Y = 32 else
"000000000000" when X = 28 AND Y = 32 else
"000000000000" when X = 29 AND Y = 32 else
"000000000000" when X = 30 AND Y = 32 else
"000000000000" when X = 31 AND Y = 32 else
"000000000000" when X = 32 AND Y = 32 else
"000000000000" when X = 33 AND Y = 32 else
"000000000000" when X = 34 AND Y = 32 else
"000000000000" when X = 35 AND Y = 32 else
"000000000000" when X = 36 AND Y = 32 else
"000000000000" when X = 37 AND Y = 32 else
"000000000000" when X = 38 AND Y = 32 else
"000000000000" when X = 39 AND Y = 32 else
"100010011101" when X = 40 AND Y = 32 else
"100010011101" when X = 41 AND Y = 32 else
"100010011101" when X = 42 AND Y = 32 else
"100010011101" when X = 43 AND Y = 32 else
"100010011101" when X = 44 AND Y = 32 else
"100010011101" when X = 45 AND Y = 32 else
"100010011101" when X = 46 AND Y = 32 else
"100010011101" when X = 47 AND Y = 32 else
"100010011101" when X = 48 AND Y = 32 else
"100010011101" when X = 49 AND Y = 32 else
"110111011111" when X = 50 AND Y = 32 else
"110111011111" when X = 51 AND Y = 32 else
"110111011111" when X = 52 AND Y = 32 else
"110111011111" when X = 53 AND Y = 32 else
"110111011111" when X = 54 AND Y = 32 else
"110111011111" when X = 55 AND Y = 32 else
"110111011111" when X = 56 AND Y = 32 else
"110111011111" when X = 57 AND Y = 32 else
"110111011111" when X = 58 AND Y = 32 else
"110111011111" when X = 59 AND Y = 32 else
"111111111111" when X = 60 AND Y = 32 else
"111111111111" when X = 61 AND Y = 32 else
"111111111111" when X = 62 AND Y = 32 else
"111111111111" when X = 63 AND Y = 32 else
"111111111111" when X = 64 AND Y = 32 else
"111111111111" when X = 65 AND Y = 32 else
"111111111111" when X = 66 AND Y = 32 else
"111111111111" when X = 67 AND Y = 32 else
"111111111111" when X = 68 AND Y = 32 else
"111111111111" when X = 69 AND Y = 32 else
"111111111111" when X = 70 AND Y = 32 else
"111111111111" when X = 71 AND Y = 32 else
"111111111111" when X = 72 AND Y = 32 else
"111111111111" when X = 73 AND Y = 32 else
"111111111111" when X = 74 AND Y = 32 else
"111111111111" when X = 75 AND Y = 32 else
"111111111111" when X = 76 AND Y = 32 else
"111111111111" when X = 77 AND Y = 32 else
"111111111111" when X = 78 AND Y = 32 else
"111111111111" when X = 79 AND Y = 32 else
"111111111111" when X = 80 AND Y = 32 else
"111111111111" when X = 81 AND Y = 32 else
"111111111111" when X = 82 AND Y = 32 else
"111111111111" when X = 83 AND Y = 32 else
"111111111111" when X = 84 AND Y = 32 else
"111111111111" when X = 85 AND Y = 32 else
"111111111111" when X = 86 AND Y = 32 else
"111111111111" when X = 87 AND Y = 32 else
"111111111111" when X = 88 AND Y = 32 else
"111111111111" when X = 89 AND Y = 32 else
"111111111111" when X = 90 AND Y = 32 else
"111111111111" when X = 91 AND Y = 32 else
"111111111111" when X = 92 AND Y = 32 else
"111111111111" when X = 93 AND Y = 32 else
"111111111111" when X = 94 AND Y = 32 else
"111111111111" when X = 95 AND Y = 32 else
"111111111111" when X = 96 AND Y = 32 else
"111111111111" when X = 97 AND Y = 32 else
"111111111111" when X = 98 AND Y = 32 else
"111111111111" when X = 99 AND Y = 32 else
"111111111111" when X = 100 AND Y = 32 else
"111111111111" when X = 101 AND Y = 32 else
"111111111111" when X = 102 AND Y = 32 else
"111111111111" when X = 103 AND Y = 32 else
"111111111111" when X = 104 AND Y = 32 else
"111111111111" when X = 105 AND Y = 32 else
"111111111111" when X = 106 AND Y = 32 else
"111111111111" when X = 107 AND Y = 32 else
"111111111111" when X = 108 AND Y = 32 else
"111111111111" when X = 109 AND Y = 32 else
"111111111111" when X = 110 AND Y = 32 else
"111111111111" when X = 111 AND Y = 32 else
"111111111111" when X = 112 AND Y = 32 else
"111111111111" when X = 113 AND Y = 32 else
"111111111111" when X = 114 AND Y = 32 else
"111111111111" when X = 115 AND Y = 32 else
"111111111111" when X = 116 AND Y = 32 else
"111111111111" when X = 117 AND Y = 32 else
"111111111111" when X = 118 AND Y = 32 else
"111111111111" when X = 119 AND Y = 32 else
"111111111111" when X = 120 AND Y = 32 else
"111111111111" when X = 121 AND Y = 32 else
"111111111111" when X = 122 AND Y = 32 else
"111111111111" when X = 123 AND Y = 32 else
"111111111111" when X = 124 AND Y = 32 else
"111111111111" when X = 125 AND Y = 32 else
"111111111111" when X = 126 AND Y = 32 else
"111111111111" when X = 127 AND Y = 32 else
"111111111111" when X = 128 AND Y = 32 else
"111111111111" when X = 129 AND Y = 32 else
"111111111111" when X = 130 AND Y = 32 else
"111111111111" when X = 131 AND Y = 32 else
"111111111111" when X = 132 AND Y = 32 else
"111111111111" when X = 133 AND Y = 32 else
"111111111111" when X = 134 AND Y = 32 else
"111111111111" when X = 135 AND Y = 32 else
"111111111111" when X = 136 AND Y = 32 else
"111111111111" when X = 137 AND Y = 32 else
"111111111111" when X = 138 AND Y = 32 else
"111111111111" when X = 139 AND Y = 32 else
"111111111111" when X = 140 AND Y = 32 else
"111111111111" when X = 141 AND Y = 32 else
"111111111111" when X = 142 AND Y = 32 else
"111111111111" when X = 143 AND Y = 32 else
"111111111111" when X = 144 AND Y = 32 else
"111111111111" when X = 145 AND Y = 32 else
"111111111111" when X = 146 AND Y = 32 else
"111111111111" when X = 147 AND Y = 32 else
"111111111111" when X = 148 AND Y = 32 else
"111111111111" when X = 149 AND Y = 32 else
"111111111111" when X = 150 AND Y = 32 else
"111111111111" when X = 151 AND Y = 32 else
"111111111111" when X = 152 AND Y = 32 else
"111111111111" when X = 153 AND Y = 32 else
"111111111111" when X = 154 AND Y = 32 else
"111111111111" when X = 155 AND Y = 32 else
"111111111111" when X = 156 AND Y = 32 else
"111111111111" when X = 157 AND Y = 32 else
"111111111111" when X = 158 AND Y = 32 else
"111111111111" when X = 159 AND Y = 32 else
"111111111111" when X = 160 AND Y = 32 else
"111111111111" when X = 161 AND Y = 32 else
"111111111111" when X = 162 AND Y = 32 else
"111111111111" when X = 163 AND Y = 32 else
"111111111111" when X = 164 AND Y = 32 else
"111111111111" when X = 165 AND Y = 32 else
"111111111111" when X = 166 AND Y = 32 else
"111111111111" when X = 167 AND Y = 32 else
"111111111111" when X = 168 AND Y = 32 else
"111111111111" when X = 169 AND Y = 32 else
"111111111111" when X = 170 AND Y = 32 else
"111111111111" when X = 171 AND Y = 32 else
"111111111111" when X = 172 AND Y = 32 else
"111111111111" when X = 173 AND Y = 32 else
"111111111111" when X = 174 AND Y = 32 else
"111111111111" when X = 175 AND Y = 32 else
"111111111111" when X = 176 AND Y = 32 else
"111111111111" when X = 177 AND Y = 32 else
"111111111111" when X = 178 AND Y = 32 else
"111111111111" when X = 179 AND Y = 32 else
"111111111111" when X = 180 AND Y = 32 else
"111111111111" when X = 181 AND Y = 32 else
"111111111111" when X = 182 AND Y = 32 else
"111111111111" when X = 183 AND Y = 32 else
"111111111111" when X = 184 AND Y = 32 else
"111111111111" when X = 185 AND Y = 32 else
"111111111111" when X = 186 AND Y = 32 else
"111111111111" when X = 187 AND Y = 32 else
"111111111111" when X = 188 AND Y = 32 else
"111111111111" when X = 189 AND Y = 32 else
"000000000000" when X = 190 AND Y = 32 else
"000000000000" when X = 191 AND Y = 32 else
"000000000000" when X = 192 AND Y = 32 else
"000000000000" when X = 193 AND Y = 32 else
"000000000000" when X = 194 AND Y = 32 else
"000000000000" when X = 195 AND Y = 32 else
"000000000000" when X = 196 AND Y = 32 else
"000000000000" when X = 197 AND Y = 32 else
"000000000000" when X = 198 AND Y = 32 else
"000000000000" when X = 199 AND Y = 32 else
"000000000000" when X = 200 AND Y = 32 else
"000000000000" when X = 201 AND Y = 32 else
"000000000000" when X = 202 AND Y = 32 else
"000000000000" when X = 203 AND Y = 32 else
"000000000000" when X = 204 AND Y = 32 else
"000000000000" when X = 205 AND Y = 32 else
"000000000000" when X = 206 AND Y = 32 else
"000000000000" when X = 207 AND Y = 32 else
"000000000000" when X = 208 AND Y = 32 else
"000000000000" when X = 209 AND Y = 32 else
"000000000000" when X = 210 AND Y = 32 else
"000000000000" when X = 211 AND Y = 32 else
"000000000000" when X = 212 AND Y = 32 else
"000000000000" when X = 213 AND Y = 32 else
"000000000000" when X = 214 AND Y = 32 else
"000000000000" when X = 215 AND Y = 32 else
"000000000000" when X = 216 AND Y = 32 else
"000000000000" when X = 217 AND Y = 32 else
"000000000000" when X = 218 AND Y = 32 else
"000000000000" when X = 219 AND Y = 32 else
"000000000000" when X = 220 AND Y = 32 else
"000000000000" when X = 221 AND Y = 32 else
"000000000000" when X = 222 AND Y = 32 else
"000000000000" when X = 223 AND Y = 32 else
"000000000000" when X = 224 AND Y = 32 else
"111111111111" when X = 225 AND Y = 32 else
"111111111111" when X = 226 AND Y = 32 else
"111111111111" when X = 227 AND Y = 32 else
"111111111111" when X = 228 AND Y = 32 else
"111111111111" when X = 229 AND Y = 32 else
"111111111111" when X = 230 AND Y = 32 else
"111111111111" when X = 231 AND Y = 32 else
"111111111111" when X = 232 AND Y = 32 else
"111111111111" when X = 233 AND Y = 32 else
"111111111111" when X = 234 AND Y = 32 else
"111111111111" when X = 235 AND Y = 32 else
"111111111111" when X = 236 AND Y = 32 else
"111111111111" when X = 237 AND Y = 32 else
"111111111111" when X = 238 AND Y = 32 else
"111111111111" when X = 239 AND Y = 32 else
"111111111111" when X = 240 AND Y = 32 else
"111111111111" when X = 241 AND Y = 32 else
"111111111111" when X = 242 AND Y = 32 else
"111111111111" when X = 243 AND Y = 32 else
"111111111111" when X = 244 AND Y = 32 else
"111111111111" when X = 245 AND Y = 32 else
"111111111111" when X = 246 AND Y = 32 else
"111111111111" when X = 247 AND Y = 32 else
"111111111111" when X = 248 AND Y = 32 else
"111111111111" when X = 249 AND Y = 32 else
"111111111111" when X = 250 AND Y = 32 else
"111111111111" when X = 251 AND Y = 32 else
"111111111111" when X = 252 AND Y = 32 else
"111111111111" when X = 253 AND Y = 32 else
"111111111111" when X = 254 AND Y = 32 else
"110111011111" when X = 255 AND Y = 32 else
"110111011111" when X = 256 AND Y = 32 else
"110111011111" when X = 257 AND Y = 32 else
"110111011111" when X = 258 AND Y = 32 else
"110111011111" when X = 259 AND Y = 32 else
"110111011111" when X = 260 AND Y = 32 else
"110111011111" when X = 261 AND Y = 32 else
"110111011111" when X = 262 AND Y = 32 else
"110111011111" when X = 263 AND Y = 32 else
"110111011111" when X = 264 AND Y = 32 else
"110111011111" when X = 265 AND Y = 32 else
"110111011111" when X = 266 AND Y = 32 else
"110111011111" when X = 267 AND Y = 32 else
"110111011111" when X = 268 AND Y = 32 else
"110111011111" when X = 269 AND Y = 32 else
"110111011111" when X = 270 AND Y = 32 else
"110111011111" when X = 271 AND Y = 32 else
"110111011111" when X = 272 AND Y = 32 else
"110111011111" when X = 273 AND Y = 32 else
"110111011111" when X = 274 AND Y = 32 else
"110111011111" when X = 275 AND Y = 32 else
"110111011111" when X = 276 AND Y = 32 else
"110111011111" when X = 277 AND Y = 32 else
"110111011111" when X = 278 AND Y = 32 else
"110111011111" when X = 279 AND Y = 32 else
"000000000000" when X = 280 AND Y = 32 else
"000000000000" when X = 281 AND Y = 32 else
"000000000000" when X = 282 AND Y = 32 else
"000000000000" when X = 283 AND Y = 32 else
"000000000000" when X = 284 AND Y = 32 else
"000000000000" when X = 285 AND Y = 32 else
"000000000000" when X = 286 AND Y = 32 else
"000000000000" when X = 287 AND Y = 32 else
"000000000000" when X = 288 AND Y = 32 else
"000000000000" when X = 289 AND Y = 32 else
"000000000000" when X = 290 AND Y = 32 else
"000000000000" when X = 291 AND Y = 32 else
"000000000000" when X = 292 AND Y = 32 else
"000000000000" when X = 293 AND Y = 32 else
"000000000000" when X = 294 AND Y = 32 else
"000000000000" when X = 295 AND Y = 32 else
"000000000000" when X = 296 AND Y = 32 else
"000000000000" when X = 297 AND Y = 32 else
"000000000000" when X = 298 AND Y = 32 else
"000000000000" when X = 299 AND Y = 32 else
"000000000000" when X = 300 AND Y = 32 else
"000000000000" when X = 301 AND Y = 32 else
"000000000000" when X = 302 AND Y = 32 else
"000000000000" when X = 303 AND Y = 32 else
"000000000000" when X = 304 AND Y = 32 else
"000000000000" when X = 305 AND Y = 32 else
"000000000000" when X = 306 AND Y = 32 else
"000000000000" when X = 307 AND Y = 32 else
"000000000000" when X = 308 AND Y = 32 else
"000000000000" when X = 309 AND Y = 32 else
"000000000000" when X = 310 AND Y = 32 else
"000000000000" when X = 311 AND Y = 32 else
"000000000000" when X = 312 AND Y = 32 else
"000000000000" when X = 313 AND Y = 32 else
"000000000000" when X = 314 AND Y = 32 else
"000000000000" when X = 315 AND Y = 32 else
"000000000000" when X = 316 AND Y = 32 else
"000000000000" when X = 317 AND Y = 32 else
"000000000000" when X = 318 AND Y = 32 else
"000000000000" when X = 319 AND Y = 32 else
"000000000000" when X = 320 AND Y = 32 else
"000000000000" when X = 321 AND Y = 32 else
"000000000000" when X = 322 AND Y = 32 else
"000000000000" when X = 323 AND Y = 32 else
"000000000000" when X = 324 AND Y = 32 else
"000000000000" when X = 0 AND Y = 33 else
"000000000000" when X = 1 AND Y = 33 else
"000000000000" when X = 2 AND Y = 33 else
"000000000000" when X = 3 AND Y = 33 else
"000000000000" when X = 4 AND Y = 33 else
"000000000000" when X = 5 AND Y = 33 else
"000000000000" when X = 6 AND Y = 33 else
"000000000000" when X = 7 AND Y = 33 else
"000000000000" when X = 8 AND Y = 33 else
"000000000000" when X = 9 AND Y = 33 else
"000000000000" when X = 10 AND Y = 33 else
"000000000000" when X = 11 AND Y = 33 else
"000000000000" when X = 12 AND Y = 33 else
"000000000000" when X = 13 AND Y = 33 else
"000000000000" when X = 14 AND Y = 33 else
"000000000000" when X = 15 AND Y = 33 else
"000000000000" when X = 16 AND Y = 33 else
"000000000000" when X = 17 AND Y = 33 else
"000000000000" when X = 18 AND Y = 33 else
"000000000000" when X = 19 AND Y = 33 else
"000000000000" when X = 20 AND Y = 33 else
"000000000000" when X = 21 AND Y = 33 else
"000000000000" when X = 22 AND Y = 33 else
"000000000000" when X = 23 AND Y = 33 else
"000000000000" when X = 24 AND Y = 33 else
"000000000000" when X = 25 AND Y = 33 else
"000000000000" when X = 26 AND Y = 33 else
"000000000000" when X = 27 AND Y = 33 else
"000000000000" when X = 28 AND Y = 33 else
"000000000000" when X = 29 AND Y = 33 else
"000000000000" when X = 30 AND Y = 33 else
"000000000000" when X = 31 AND Y = 33 else
"000000000000" when X = 32 AND Y = 33 else
"000000000000" when X = 33 AND Y = 33 else
"000000000000" when X = 34 AND Y = 33 else
"000000000000" when X = 35 AND Y = 33 else
"000000000000" when X = 36 AND Y = 33 else
"000000000000" when X = 37 AND Y = 33 else
"000000000000" when X = 38 AND Y = 33 else
"000000000000" when X = 39 AND Y = 33 else
"100010011101" when X = 40 AND Y = 33 else
"100010011101" when X = 41 AND Y = 33 else
"100010011101" when X = 42 AND Y = 33 else
"100010011101" when X = 43 AND Y = 33 else
"100010011101" when X = 44 AND Y = 33 else
"100010011101" when X = 45 AND Y = 33 else
"100010011101" when X = 46 AND Y = 33 else
"100010011101" when X = 47 AND Y = 33 else
"100010011101" when X = 48 AND Y = 33 else
"100010011101" when X = 49 AND Y = 33 else
"110111011111" when X = 50 AND Y = 33 else
"110111011111" when X = 51 AND Y = 33 else
"110111011111" when X = 52 AND Y = 33 else
"110111011111" when X = 53 AND Y = 33 else
"110111011111" when X = 54 AND Y = 33 else
"110111011111" when X = 55 AND Y = 33 else
"110111011111" when X = 56 AND Y = 33 else
"110111011111" when X = 57 AND Y = 33 else
"110111011111" when X = 58 AND Y = 33 else
"110111011111" when X = 59 AND Y = 33 else
"111111111111" when X = 60 AND Y = 33 else
"111111111111" when X = 61 AND Y = 33 else
"111111111111" when X = 62 AND Y = 33 else
"111111111111" when X = 63 AND Y = 33 else
"111111111111" when X = 64 AND Y = 33 else
"111111111111" when X = 65 AND Y = 33 else
"111111111111" when X = 66 AND Y = 33 else
"111111111111" when X = 67 AND Y = 33 else
"111111111111" when X = 68 AND Y = 33 else
"111111111111" when X = 69 AND Y = 33 else
"111111111111" when X = 70 AND Y = 33 else
"111111111111" when X = 71 AND Y = 33 else
"111111111111" when X = 72 AND Y = 33 else
"111111111111" when X = 73 AND Y = 33 else
"111111111111" when X = 74 AND Y = 33 else
"111111111111" when X = 75 AND Y = 33 else
"111111111111" when X = 76 AND Y = 33 else
"111111111111" when X = 77 AND Y = 33 else
"111111111111" when X = 78 AND Y = 33 else
"111111111111" when X = 79 AND Y = 33 else
"111111111111" when X = 80 AND Y = 33 else
"111111111111" when X = 81 AND Y = 33 else
"111111111111" when X = 82 AND Y = 33 else
"111111111111" when X = 83 AND Y = 33 else
"111111111111" when X = 84 AND Y = 33 else
"111111111111" when X = 85 AND Y = 33 else
"111111111111" when X = 86 AND Y = 33 else
"111111111111" when X = 87 AND Y = 33 else
"111111111111" when X = 88 AND Y = 33 else
"111111111111" when X = 89 AND Y = 33 else
"111111111111" when X = 90 AND Y = 33 else
"111111111111" when X = 91 AND Y = 33 else
"111111111111" when X = 92 AND Y = 33 else
"111111111111" when X = 93 AND Y = 33 else
"111111111111" when X = 94 AND Y = 33 else
"111111111111" when X = 95 AND Y = 33 else
"111111111111" when X = 96 AND Y = 33 else
"111111111111" when X = 97 AND Y = 33 else
"111111111111" when X = 98 AND Y = 33 else
"111111111111" when X = 99 AND Y = 33 else
"111111111111" when X = 100 AND Y = 33 else
"111111111111" when X = 101 AND Y = 33 else
"111111111111" when X = 102 AND Y = 33 else
"111111111111" when X = 103 AND Y = 33 else
"111111111111" when X = 104 AND Y = 33 else
"111111111111" when X = 105 AND Y = 33 else
"111111111111" when X = 106 AND Y = 33 else
"111111111111" when X = 107 AND Y = 33 else
"111111111111" when X = 108 AND Y = 33 else
"111111111111" when X = 109 AND Y = 33 else
"111111111111" when X = 110 AND Y = 33 else
"111111111111" when X = 111 AND Y = 33 else
"111111111111" when X = 112 AND Y = 33 else
"111111111111" when X = 113 AND Y = 33 else
"111111111111" when X = 114 AND Y = 33 else
"111111111111" when X = 115 AND Y = 33 else
"111111111111" when X = 116 AND Y = 33 else
"111111111111" when X = 117 AND Y = 33 else
"111111111111" when X = 118 AND Y = 33 else
"111111111111" when X = 119 AND Y = 33 else
"111111111111" when X = 120 AND Y = 33 else
"111111111111" when X = 121 AND Y = 33 else
"111111111111" when X = 122 AND Y = 33 else
"111111111111" when X = 123 AND Y = 33 else
"111111111111" when X = 124 AND Y = 33 else
"111111111111" when X = 125 AND Y = 33 else
"111111111111" when X = 126 AND Y = 33 else
"111111111111" when X = 127 AND Y = 33 else
"111111111111" when X = 128 AND Y = 33 else
"111111111111" when X = 129 AND Y = 33 else
"111111111111" when X = 130 AND Y = 33 else
"111111111111" when X = 131 AND Y = 33 else
"111111111111" when X = 132 AND Y = 33 else
"111111111111" when X = 133 AND Y = 33 else
"111111111111" when X = 134 AND Y = 33 else
"111111111111" when X = 135 AND Y = 33 else
"111111111111" when X = 136 AND Y = 33 else
"111111111111" when X = 137 AND Y = 33 else
"111111111111" when X = 138 AND Y = 33 else
"111111111111" when X = 139 AND Y = 33 else
"111111111111" when X = 140 AND Y = 33 else
"111111111111" when X = 141 AND Y = 33 else
"111111111111" when X = 142 AND Y = 33 else
"111111111111" when X = 143 AND Y = 33 else
"111111111111" when X = 144 AND Y = 33 else
"111111111111" when X = 145 AND Y = 33 else
"111111111111" when X = 146 AND Y = 33 else
"111111111111" when X = 147 AND Y = 33 else
"111111111111" when X = 148 AND Y = 33 else
"111111111111" when X = 149 AND Y = 33 else
"111111111111" when X = 150 AND Y = 33 else
"111111111111" when X = 151 AND Y = 33 else
"111111111111" when X = 152 AND Y = 33 else
"111111111111" when X = 153 AND Y = 33 else
"111111111111" when X = 154 AND Y = 33 else
"111111111111" when X = 155 AND Y = 33 else
"111111111111" when X = 156 AND Y = 33 else
"111111111111" when X = 157 AND Y = 33 else
"111111111111" when X = 158 AND Y = 33 else
"111111111111" when X = 159 AND Y = 33 else
"111111111111" when X = 160 AND Y = 33 else
"111111111111" when X = 161 AND Y = 33 else
"111111111111" when X = 162 AND Y = 33 else
"111111111111" when X = 163 AND Y = 33 else
"111111111111" when X = 164 AND Y = 33 else
"111111111111" when X = 165 AND Y = 33 else
"111111111111" when X = 166 AND Y = 33 else
"111111111111" when X = 167 AND Y = 33 else
"111111111111" when X = 168 AND Y = 33 else
"111111111111" when X = 169 AND Y = 33 else
"111111111111" when X = 170 AND Y = 33 else
"111111111111" when X = 171 AND Y = 33 else
"111111111111" when X = 172 AND Y = 33 else
"111111111111" when X = 173 AND Y = 33 else
"111111111111" when X = 174 AND Y = 33 else
"111111111111" when X = 175 AND Y = 33 else
"111111111111" when X = 176 AND Y = 33 else
"111111111111" when X = 177 AND Y = 33 else
"111111111111" when X = 178 AND Y = 33 else
"111111111111" when X = 179 AND Y = 33 else
"111111111111" when X = 180 AND Y = 33 else
"111111111111" when X = 181 AND Y = 33 else
"111111111111" when X = 182 AND Y = 33 else
"111111111111" when X = 183 AND Y = 33 else
"111111111111" when X = 184 AND Y = 33 else
"111111111111" when X = 185 AND Y = 33 else
"111111111111" when X = 186 AND Y = 33 else
"111111111111" when X = 187 AND Y = 33 else
"111111111111" when X = 188 AND Y = 33 else
"111111111111" when X = 189 AND Y = 33 else
"000000000000" when X = 190 AND Y = 33 else
"000000000000" when X = 191 AND Y = 33 else
"000000000000" when X = 192 AND Y = 33 else
"000000000000" when X = 193 AND Y = 33 else
"000000000000" when X = 194 AND Y = 33 else
"000000000000" when X = 195 AND Y = 33 else
"000000000000" when X = 196 AND Y = 33 else
"000000000000" when X = 197 AND Y = 33 else
"000000000000" when X = 198 AND Y = 33 else
"000000000000" when X = 199 AND Y = 33 else
"000000000000" when X = 200 AND Y = 33 else
"000000000000" when X = 201 AND Y = 33 else
"000000000000" when X = 202 AND Y = 33 else
"000000000000" when X = 203 AND Y = 33 else
"000000000000" when X = 204 AND Y = 33 else
"000000000000" when X = 205 AND Y = 33 else
"000000000000" when X = 206 AND Y = 33 else
"000000000000" when X = 207 AND Y = 33 else
"000000000000" when X = 208 AND Y = 33 else
"000000000000" when X = 209 AND Y = 33 else
"000000000000" when X = 210 AND Y = 33 else
"000000000000" when X = 211 AND Y = 33 else
"000000000000" when X = 212 AND Y = 33 else
"000000000000" when X = 213 AND Y = 33 else
"000000000000" when X = 214 AND Y = 33 else
"000000000000" when X = 215 AND Y = 33 else
"000000000000" when X = 216 AND Y = 33 else
"000000000000" when X = 217 AND Y = 33 else
"000000000000" when X = 218 AND Y = 33 else
"000000000000" when X = 219 AND Y = 33 else
"000000000000" when X = 220 AND Y = 33 else
"000000000000" when X = 221 AND Y = 33 else
"000000000000" when X = 222 AND Y = 33 else
"000000000000" when X = 223 AND Y = 33 else
"000000000000" when X = 224 AND Y = 33 else
"111111111111" when X = 225 AND Y = 33 else
"111111111111" when X = 226 AND Y = 33 else
"111111111111" when X = 227 AND Y = 33 else
"111111111111" when X = 228 AND Y = 33 else
"111111111111" when X = 229 AND Y = 33 else
"111111111111" when X = 230 AND Y = 33 else
"111111111111" when X = 231 AND Y = 33 else
"111111111111" when X = 232 AND Y = 33 else
"111111111111" when X = 233 AND Y = 33 else
"111111111111" when X = 234 AND Y = 33 else
"111111111111" when X = 235 AND Y = 33 else
"111111111111" when X = 236 AND Y = 33 else
"111111111111" when X = 237 AND Y = 33 else
"111111111111" when X = 238 AND Y = 33 else
"111111111111" when X = 239 AND Y = 33 else
"111111111111" when X = 240 AND Y = 33 else
"111111111111" when X = 241 AND Y = 33 else
"111111111111" when X = 242 AND Y = 33 else
"111111111111" when X = 243 AND Y = 33 else
"111111111111" when X = 244 AND Y = 33 else
"111111111111" when X = 245 AND Y = 33 else
"111111111111" when X = 246 AND Y = 33 else
"111111111111" when X = 247 AND Y = 33 else
"111111111111" when X = 248 AND Y = 33 else
"111111111111" when X = 249 AND Y = 33 else
"111111111111" when X = 250 AND Y = 33 else
"111111111111" when X = 251 AND Y = 33 else
"111111111111" when X = 252 AND Y = 33 else
"111111111111" when X = 253 AND Y = 33 else
"111111111111" when X = 254 AND Y = 33 else
"110111011111" when X = 255 AND Y = 33 else
"110111011111" when X = 256 AND Y = 33 else
"110111011111" when X = 257 AND Y = 33 else
"110111011111" when X = 258 AND Y = 33 else
"110111011111" when X = 259 AND Y = 33 else
"110111011111" when X = 260 AND Y = 33 else
"110111011111" when X = 261 AND Y = 33 else
"110111011111" when X = 262 AND Y = 33 else
"110111011111" when X = 263 AND Y = 33 else
"110111011111" when X = 264 AND Y = 33 else
"110111011111" when X = 265 AND Y = 33 else
"110111011111" when X = 266 AND Y = 33 else
"110111011111" when X = 267 AND Y = 33 else
"110111011111" when X = 268 AND Y = 33 else
"110111011111" when X = 269 AND Y = 33 else
"110111011111" when X = 270 AND Y = 33 else
"110111011111" when X = 271 AND Y = 33 else
"110111011111" when X = 272 AND Y = 33 else
"110111011111" when X = 273 AND Y = 33 else
"110111011111" when X = 274 AND Y = 33 else
"110111011111" when X = 275 AND Y = 33 else
"110111011111" when X = 276 AND Y = 33 else
"110111011111" when X = 277 AND Y = 33 else
"110111011111" when X = 278 AND Y = 33 else
"110111011111" when X = 279 AND Y = 33 else
"000000000000" when X = 280 AND Y = 33 else
"000000000000" when X = 281 AND Y = 33 else
"000000000000" when X = 282 AND Y = 33 else
"000000000000" when X = 283 AND Y = 33 else
"000000000000" when X = 284 AND Y = 33 else
"000000000000" when X = 285 AND Y = 33 else
"000000000000" when X = 286 AND Y = 33 else
"000000000000" when X = 287 AND Y = 33 else
"000000000000" when X = 288 AND Y = 33 else
"000000000000" when X = 289 AND Y = 33 else
"000000000000" when X = 290 AND Y = 33 else
"000000000000" when X = 291 AND Y = 33 else
"000000000000" when X = 292 AND Y = 33 else
"000000000000" when X = 293 AND Y = 33 else
"000000000000" when X = 294 AND Y = 33 else
"000000000000" when X = 295 AND Y = 33 else
"000000000000" when X = 296 AND Y = 33 else
"000000000000" when X = 297 AND Y = 33 else
"000000000000" when X = 298 AND Y = 33 else
"000000000000" when X = 299 AND Y = 33 else
"000000000000" when X = 300 AND Y = 33 else
"000000000000" when X = 301 AND Y = 33 else
"000000000000" when X = 302 AND Y = 33 else
"000000000000" when X = 303 AND Y = 33 else
"000000000000" when X = 304 AND Y = 33 else
"000000000000" when X = 305 AND Y = 33 else
"000000000000" when X = 306 AND Y = 33 else
"000000000000" when X = 307 AND Y = 33 else
"000000000000" when X = 308 AND Y = 33 else
"000000000000" when X = 309 AND Y = 33 else
"000000000000" when X = 310 AND Y = 33 else
"000000000000" when X = 311 AND Y = 33 else
"000000000000" when X = 312 AND Y = 33 else
"000000000000" when X = 313 AND Y = 33 else
"000000000000" when X = 314 AND Y = 33 else
"000000000000" when X = 315 AND Y = 33 else
"000000000000" when X = 316 AND Y = 33 else
"000000000000" when X = 317 AND Y = 33 else
"000000000000" when X = 318 AND Y = 33 else
"000000000000" when X = 319 AND Y = 33 else
"000000000000" when X = 320 AND Y = 33 else
"000000000000" when X = 321 AND Y = 33 else
"000000000000" when X = 322 AND Y = 33 else
"000000000000" when X = 323 AND Y = 33 else
"000000000000" when X = 324 AND Y = 33 else
"000000000000" when X = 0 AND Y = 34 else
"000000000000" when X = 1 AND Y = 34 else
"000000000000" when X = 2 AND Y = 34 else
"000000000000" when X = 3 AND Y = 34 else
"000000000000" when X = 4 AND Y = 34 else
"000000000000" when X = 5 AND Y = 34 else
"000000000000" when X = 6 AND Y = 34 else
"000000000000" when X = 7 AND Y = 34 else
"000000000000" when X = 8 AND Y = 34 else
"000000000000" when X = 9 AND Y = 34 else
"000000000000" when X = 10 AND Y = 34 else
"000000000000" when X = 11 AND Y = 34 else
"000000000000" when X = 12 AND Y = 34 else
"000000000000" when X = 13 AND Y = 34 else
"000000000000" when X = 14 AND Y = 34 else
"000000000000" when X = 15 AND Y = 34 else
"000000000000" when X = 16 AND Y = 34 else
"000000000000" when X = 17 AND Y = 34 else
"000000000000" when X = 18 AND Y = 34 else
"000000000000" when X = 19 AND Y = 34 else
"000000000000" when X = 20 AND Y = 34 else
"000000000000" when X = 21 AND Y = 34 else
"000000000000" when X = 22 AND Y = 34 else
"000000000000" when X = 23 AND Y = 34 else
"000000000000" when X = 24 AND Y = 34 else
"000000000000" when X = 25 AND Y = 34 else
"000000000000" when X = 26 AND Y = 34 else
"000000000000" when X = 27 AND Y = 34 else
"000000000000" when X = 28 AND Y = 34 else
"000000000000" when X = 29 AND Y = 34 else
"000000000000" when X = 30 AND Y = 34 else
"000000000000" when X = 31 AND Y = 34 else
"000000000000" when X = 32 AND Y = 34 else
"000000000000" when X = 33 AND Y = 34 else
"000000000000" when X = 34 AND Y = 34 else
"000000000000" when X = 35 AND Y = 34 else
"000000000000" when X = 36 AND Y = 34 else
"000000000000" when X = 37 AND Y = 34 else
"000000000000" when X = 38 AND Y = 34 else
"000000000000" when X = 39 AND Y = 34 else
"100010011101" when X = 40 AND Y = 34 else
"100010011101" when X = 41 AND Y = 34 else
"100010011101" when X = 42 AND Y = 34 else
"100010011101" when X = 43 AND Y = 34 else
"100010011101" when X = 44 AND Y = 34 else
"100010011101" when X = 45 AND Y = 34 else
"100010011101" when X = 46 AND Y = 34 else
"100010011101" when X = 47 AND Y = 34 else
"100010011101" when X = 48 AND Y = 34 else
"100010011101" when X = 49 AND Y = 34 else
"110111011111" when X = 50 AND Y = 34 else
"110111011111" when X = 51 AND Y = 34 else
"110111011111" when X = 52 AND Y = 34 else
"110111011111" when X = 53 AND Y = 34 else
"110111011111" when X = 54 AND Y = 34 else
"110111011111" when X = 55 AND Y = 34 else
"110111011111" when X = 56 AND Y = 34 else
"110111011111" when X = 57 AND Y = 34 else
"110111011111" when X = 58 AND Y = 34 else
"110111011111" when X = 59 AND Y = 34 else
"111111111111" when X = 60 AND Y = 34 else
"111111111111" when X = 61 AND Y = 34 else
"111111111111" when X = 62 AND Y = 34 else
"111111111111" when X = 63 AND Y = 34 else
"111111111111" when X = 64 AND Y = 34 else
"111111111111" when X = 65 AND Y = 34 else
"111111111111" when X = 66 AND Y = 34 else
"111111111111" when X = 67 AND Y = 34 else
"111111111111" when X = 68 AND Y = 34 else
"111111111111" when X = 69 AND Y = 34 else
"111111111111" when X = 70 AND Y = 34 else
"111111111111" when X = 71 AND Y = 34 else
"111111111111" when X = 72 AND Y = 34 else
"111111111111" when X = 73 AND Y = 34 else
"111111111111" when X = 74 AND Y = 34 else
"111111111111" when X = 75 AND Y = 34 else
"111111111111" when X = 76 AND Y = 34 else
"111111111111" when X = 77 AND Y = 34 else
"111111111111" when X = 78 AND Y = 34 else
"111111111111" when X = 79 AND Y = 34 else
"111111111111" when X = 80 AND Y = 34 else
"111111111111" when X = 81 AND Y = 34 else
"111111111111" when X = 82 AND Y = 34 else
"111111111111" when X = 83 AND Y = 34 else
"111111111111" when X = 84 AND Y = 34 else
"111111111111" when X = 85 AND Y = 34 else
"111111111111" when X = 86 AND Y = 34 else
"111111111111" when X = 87 AND Y = 34 else
"111111111111" when X = 88 AND Y = 34 else
"111111111111" when X = 89 AND Y = 34 else
"111111111111" when X = 90 AND Y = 34 else
"111111111111" when X = 91 AND Y = 34 else
"111111111111" when X = 92 AND Y = 34 else
"111111111111" when X = 93 AND Y = 34 else
"111111111111" when X = 94 AND Y = 34 else
"111111111111" when X = 95 AND Y = 34 else
"111111111111" when X = 96 AND Y = 34 else
"111111111111" when X = 97 AND Y = 34 else
"111111111111" when X = 98 AND Y = 34 else
"111111111111" when X = 99 AND Y = 34 else
"111111111111" when X = 100 AND Y = 34 else
"111111111111" when X = 101 AND Y = 34 else
"111111111111" when X = 102 AND Y = 34 else
"111111111111" when X = 103 AND Y = 34 else
"111111111111" when X = 104 AND Y = 34 else
"111111111111" when X = 105 AND Y = 34 else
"111111111111" when X = 106 AND Y = 34 else
"111111111111" when X = 107 AND Y = 34 else
"111111111111" when X = 108 AND Y = 34 else
"111111111111" when X = 109 AND Y = 34 else
"111111111111" when X = 110 AND Y = 34 else
"111111111111" when X = 111 AND Y = 34 else
"111111111111" when X = 112 AND Y = 34 else
"111111111111" when X = 113 AND Y = 34 else
"111111111111" when X = 114 AND Y = 34 else
"111111111111" when X = 115 AND Y = 34 else
"111111111111" when X = 116 AND Y = 34 else
"111111111111" when X = 117 AND Y = 34 else
"111111111111" when X = 118 AND Y = 34 else
"111111111111" when X = 119 AND Y = 34 else
"111111111111" when X = 120 AND Y = 34 else
"111111111111" when X = 121 AND Y = 34 else
"111111111111" when X = 122 AND Y = 34 else
"111111111111" when X = 123 AND Y = 34 else
"111111111111" when X = 124 AND Y = 34 else
"111111111111" when X = 125 AND Y = 34 else
"111111111111" when X = 126 AND Y = 34 else
"111111111111" when X = 127 AND Y = 34 else
"111111111111" when X = 128 AND Y = 34 else
"111111111111" when X = 129 AND Y = 34 else
"111111111111" when X = 130 AND Y = 34 else
"111111111111" when X = 131 AND Y = 34 else
"111111111111" when X = 132 AND Y = 34 else
"111111111111" when X = 133 AND Y = 34 else
"111111111111" when X = 134 AND Y = 34 else
"111111111111" when X = 135 AND Y = 34 else
"111111111111" when X = 136 AND Y = 34 else
"111111111111" when X = 137 AND Y = 34 else
"111111111111" when X = 138 AND Y = 34 else
"111111111111" when X = 139 AND Y = 34 else
"111111111111" when X = 140 AND Y = 34 else
"111111111111" when X = 141 AND Y = 34 else
"111111111111" when X = 142 AND Y = 34 else
"111111111111" when X = 143 AND Y = 34 else
"111111111111" when X = 144 AND Y = 34 else
"111111111111" when X = 145 AND Y = 34 else
"111111111111" when X = 146 AND Y = 34 else
"111111111111" when X = 147 AND Y = 34 else
"111111111111" when X = 148 AND Y = 34 else
"111111111111" when X = 149 AND Y = 34 else
"111111111111" when X = 150 AND Y = 34 else
"111111111111" when X = 151 AND Y = 34 else
"111111111111" when X = 152 AND Y = 34 else
"111111111111" when X = 153 AND Y = 34 else
"111111111111" when X = 154 AND Y = 34 else
"111111111111" when X = 155 AND Y = 34 else
"111111111111" when X = 156 AND Y = 34 else
"111111111111" when X = 157 AND Y = 34 else
"111111111111" when X = 158 AND Y = 34 else
"111111111111" when X = 159 AND Y = 34 else
"111111111111" when X = 160 AND Y = 34 else
"111111111111" when X = 161 AND Y = 34 else
"111111111111" when X = 162 AND Y = 34 else
"111111111111" when X = 163 AND Y = 34 else
"111111111111" when X = 164 AND Y = 34 else
"111111111111" when X = 165 AND Y = 34 else
"111111111111" when X = 166 AND Y = 34 else
"111111111111" when X = 167 AND Y = 34 else
"111111111111" when X = 168 AND Y = 34 else
"111111111111" when X = 169 AND Y = 34 else
"111111111111" when X = 170 AND Y = 34 else
"111111111111" when X = 171 AND Y = 34 else
"111111111111" when X = 172 AND Y = 34 else
"111111111111" when X = 173 AND Y = 34 else
"111111111111" when X = 174 AND Y = 34 else
"111111111111" when X = 175 AND Y = 34 else
"111111111111" when X = 176 AND Y = 34 else
"111111111111" when X = 177 AND Y = 34 else
"111111111111" when X = 178 AND Y = 34 else
"111111111111" when X = 179 AND Y = 34 else
"111111111111" when X = 180 AND Y = 34 else
"111111111111" when X = 181 AND Y = 34 else
"111111111111" when X = 182 AND Y = 34 else
"111111111111" when X = 183 AND Y = 34 else
"111111111111" when X = 184 AND Y = 34 else
"111111111111" when X = 185 AND Y = 34 else
"111111111111" when X = 186 AND Y = 34 else
"111111111111" when X = 187 AND Y = 34 else
"111111111111" when X = 188 AND Y = 34 else
"111111111111" when X = 189 AND Y = 34 else
"000000000000" when X = 190 AND Y = 34 else
"000000000000" when X = 191 AND Y = 34 else
"000000000000" when X = 192 AND Y = 34 else
"000000000000" when X = 193 AND Y = 34 else
"000000000000" when X = 194 AND Y = 34 else
"000000000000" when X = 195 AND Y = 34 else
"000000000000" when X = 196 AND Y = 34 else
"000000000000" when X = 197 AND Y = 34 else
"000000000000" when X = 198 AND Y = 34 else
"000000000000" when X = 199 AND Y = 34 else
"000000000000" when X = 200 AND Y = 34 else
"000000000000" when X = 201 AND Y = 34 else
"000000000000" when X = 202 AND Y = 34 else
"000000000000" when X = 203 AND Y = 34 else
"000000000000" when X = 204 AND Y = 34 else
"000000000000" when X = 205 AND Y = 34 else
"000000000000" when X = 206 AND Y = 34 else
"000000000000" when X = 207 AND Y = 34 else
"000000000000" when X = 208 AND Y = 34 else
"000000000000" when X = 209 AND Y = 34 else
"000000000000" when X = 210 AND Y = 34 else
"000000000000" when X = 211 AND Y = 34 else
"000000000000" when X = 212 AND Y = 34 else
"000000000000" when X = 213 AND Y = 34 else
"000000000000" when X = 214 AND Y = 34 else
"000000000000" when X = 215 AND Y = 34 else
"000000000000" when X = 216 AND Y = 34 else
"000000000000" when X = 217 AND Y = 34 else
"000000000000" when X = 218 AND Y = 34 else
"000000000000" when X = 219 AND Y = 34 else
"000000000000" when X = 220 AND Y = 34 else
"000000000000" when X = 221 AND Y = 34 else
"000000000000" when X = 222 AND Y = 34 else
"000000000000" when X = 223 AND Y = 34 else
"000000000000" when X = 224 AND Y = 34 else
"111111111111" when X = 225 AND Y = 34 else
"111111111111" when X = 226 AND Y = 34 else
"111111111111" when X = 227 AND Y = 34 else
"111111111111" when X = 228 AND Y = 34 else
"111111111111" when X = 229 AND Y = 34 else
"111111111111" when X = 230 AND Y = 34 else
"111111111111" when X = 231 AND Y = 34 else
"111111111111" when X = 232 AND Y = 34 else
"111111111111" when X = 233 AND Y = 34 else
"111111111111" when X = 234 AND Y = 34 else
"111111111111" when X = 235 AND Y = 34 else
"111111111111" when X = 236 AND Y = 34 else
"111111111111" when X = 237 AND Y = 34 else
"111111111111" when X = 238 AND Y = 34 else
"111111111111" when X = 239 AND Y = 34 else
"111111111111" when X = 240 AND Y = 34 else
"111111111111" when X = 241 AND Y = 34 else
"111111111111" when X = 242 AND Y = 34 else
"111111111111" when X = 243 AND Y = 34 else
"111111111111" when X = 244 AND Y = 34 else
"111111111111" when X = 245 AND Y = 34 else
"111111111111" when X = 246 AND Y = 34 else
"111111111111" when X = 247 AND Y = 34 else
"111111111111" when X = 248 AND Y = 34 else
"111111111111" when X = 249 AND Y = 34 else
"111111111111" when X = 250 AND Y = 34 else
"111111111111" when X = 251 AND Y = 34 else
"111111111111" when X = 252 AND Y = 34 else
"111111111111" when X = 253 AND Y = 34 else
"111111111111" when X = 254 AND Y = 34 else
"110111011111" when X = 255 AND Y = 34 else
"110111011111" when X = 256 AND Y = 34 else
"110111011111" when X = 257 AND Y = 34 else
"110111011111" when X = 258 AND Y = 34 else
"110111011111" when X = 259 AND Y = 34 else
"110111011111" when X = 260 AND Y = 34 else
"110111011111" when X = 261 AND Y = 34 else
"110111011111" when X = 262 AND Y = 34 else
"110111011111" when X = 263 AND Y = 34 else
"110111011111" when X = 264 AND Y = 34 else
"110111011111" when X = 265 AND Y = 34 else
"110111011111" when X = 266 AND Y = 34 else
"110111011111" when X = 267 AND Y = 34 else
"110111011111" when X = 268 AND Y = 34 else
"110111011111" when X = 269 AND Y = 34 else
"110111011111" when X = 270 AND Y = 34 else
"110111011111" when X = 271 AND Y = 34 else
"110111011111" when X = 272 AND Y = 34 else
"110111011111" when X = 273 AND Y = 34 else
"110111011111" when X = 274 AND Y = 34 else
"110111011111" when X = 275 AND Y = 34 else
"110111011111" when X = 276 AND Y = 34 else
"110111011111" when X = 277 AND Y = 34 else
"110111011111" when X = 278 AND Y = 34 else
"110111011111" when X = 279 AND Y = 34 else
"000000000000" when X = 280 AND Y = 34 else
"000000000000" when X = 281 AND Y = 34 else
"000000000000" when X = 282 AND Y = 34 else
"000000000000" when X = 283 AND Y = 34 else
"000000000000" when X = 284 AND Y = 34 else
"000000000000" when X = 285 AND Y = 34 else
"000000000000" when X = 286 AND Y = 34 else
"000000000000" when X = 287 AND Y = 34 else
"000000000000" when X = 288 AND Y = 34 else
"000000000000" when X = 289 AND Y = 34 else
"000000000000" when X = 290 AND Y = 34 else
"000000000000" when X = 291 AND Y = 34 else
"000000000000" when X = 292 AND Y = 34 else
"000000000000" when X = 293 AND Y = 34 else
"000000000000" when X = 294 AND Y = 34 else
"000000000000" when X = 295 AND Y = 34 else
"000000000000" when X = 296 AND Y = 34 else
"000000000000" when X = 297 AND Y = 34 else
"000000000000" when X = 298 AND Y = 34 else
"000000000000" when X = 299 AND Y = 34 else
"000000000000" when X = 300 AND Y = 34 else
"000000000000" when X = 301 AND Y = 34 else
"000000000000" when X = 302 AND Y = 34 else
"000000000000" when X = 303 AND Y = 34 else
"000000000000" when X = 304 AND Y = 34 else
"000000000000" when X = 305 AND Y = 34 else
"000000000000" when X = 306 AND Y = 34 else
"000000000000" when X = 307 AND Y = 34 else
"000000000000" when X = 308 AND Y = 34 else
"000000000000" when X = 309 AND Y = 34 else
"000000000000" when X = 310 AND Y = 34 else
"000000000000" when X = 311 AND Y = 34 else
"000000000000" when X = 312 AND Y = 34 else
"000000000000" when X = 313 AND Y = 34 else
"000000000000" when X = 314 AND Y = 34 else
"000000000000" when X = 315 AND Y = 34 else
"000000000000" when X = 316 AND Y = 34 else
"000000000000" when X = 317 AND Y = 34 else
"000000000000" when X = 318 AND Y = 34 else
"000000000000" when X = 319 AND Y = 34 else
"000000000000" when X = 320 AND Y = 34 else
"000000000000" when X = 321 AND Y = 34 else
"000000000000" when X = 322 AND Y = 34 else
"000000000000" when X = 323 AND Y = 34 else
"000000000000" when X = 324 AND Y = 34 else
"000000000000" when X = 0 AND Y = 35 else
"000000000000" when X = 1 AND Y = 35 else
"000000000000" when X = 2 AND Y = 35 else
"000000000000" when X = 3 AND Y = 35 else
"000000000000" when X = 4 AND Y = 35 else
"000000000000" when X = 5 AND Y = 35 else
"000000000000" when X = 6 AND Y = 35 else
"000000000000" when X = 7 AND Y = 35 else
"000000000000" when X = 8 AND Y = 35 else
"000000000000" when X = 9 AND Y = 35 else
"000000000000" when X = 10 AND Y = 35 else
"000000000000" when X = 11 AND Y = 35 else
"000000000000" when X = 12 AND Y = 35 else
"000000000000" when X = 13 AND Y = 35 else
"000000000000" when X = 14 AND Y = 35 else
"000000000000" when X = 15 AND Y = 35 else
"000000000000" when X = 16 AND Y = 35 else
"000000000000" when X = 17 AND Y = 35 else
"000000000000" when X = 18 AND Y = 35 else
"000000000000" when X = 19 AND Y = 35 else
"000000000000" when X = 20 AND Y = 35 else
"000000000000" when X = 21 AND Y = 35 else
"000000000000" when X = 22 AND Y = 35 else
"000000000000" when X = 23 AND Y = 35 else
"000000000000" when X = 24 AND Y = 35 else
"000000000000" when X = 25 AND Y = 35 else
"000000000000" when X = 26 AND Y = 35 else
"000000000000" when X = 27 AND Y = 35 else
"000000000000" when X = 28 AND Y = 35 else
"000000000000" when X = 29 AND Y = 35 else
"000000000000" when X = 30 AND Y = 35 else
"000000000000" when X = 31 AND Y = 35 else
"000000000000" when X = 32 AND Y = 35 else
"000000000000" when X = 33 AND Y = 35 else
"000000000000" when X = 34 AND Y = 35 else
"000000000000" when X = 35 AND Y = 35 else
"000000000000" when X = 36 AND Y = 35 else
"000000000000" when X = 37 AND Y = 35 else
"000000000000" when X = 38 AND Y = 35 else
"000000000000" when X = 39 AND Y = 35 else
"100010011101" when X = 40 AND Y = 35 else
"100010011101" when X = 41 AND Y = 35 else
"100010011101" when X = 42 AND Y = 35 else
"100010011101" when X = 43 AND Y = 35 else
"100010011101" when X = 44 AND Y = 35 else
"100010011101" when X = 45 AND Y = 35 else
"100010011101" when X = 46 AND Y = 35 else
"100010011101" when X = 47 AND Y = 35 else
"100010011101" when X = 48 AND Y = 35 else
"100010011101" when X = 49 AND Y = 35 else
"110111011111" when X = 50 AND Y = 35 else
"110111011111" when X = 51 AND Y = 35 else
"110111011111" when X = 52 AND Y = 35 else
"110111011111" when X = 53 AND Y = 35 else
"110111011111" when X = 54 AND Y = 35 else
"110111011111" when X = 55 AND Y = 35 else
"110111011111" when X = 56 AND Y = 35 else
"110111011111" when X = 57 AND Y = 35 else
"110111011111" when X = 58 AND Y = 35 else
"110111011111" when X = 59 AND Y = 35 else
"111111111111" when X = 60 AND Y = 35 else
"111111111111" when X = 61 AND Y = 35 else
"111111111111" when X = 62 AND Y = 35 else
"111111111111" when X = 63 AND Y = 35 else
"111111111111" when X = 64 AND Y = 35 else
"111111111111" when X = 65 AND Y = 35 else
"111111111111" when X = 66 AND Y = 35 else
"111111111111" when X = 67 AND Y = 35 else
"111111111111" when X = 68 AND Y = 35 else
"111111111111" when X = 69 AND Y = 35 else
"111111111111" when X = 70 AND Y = 35 else
"111111111111" when X = 71 AND Y = 35 else
"111111111111" when X = 72 AND Y = 35 else
"111111111111" when X = 73 AND Y = 35 else
"111111111111" when X = 74 AND Y = 35 else
"111111111111" when X = 75 AND Y = 35 else
"111111111111" when X = 76 AND Y = 35 else
"111111111111" when X = 77 AND Y = 35 else
"111111111111" when X = 78 AND Y = 35 else
"111111111111" when X = 79 AND Y = 35 else
"111111111111" when X = 80 AND Y = 35 else
"111111111111" when X = 81 AND Y = 35 else
"111111111111" when X = 82 AND Y = 35 else
"111111111111" when X = 83 AND Y = 35 else
"111111111111" when X = 84 AND Y = 35 else
"111111111111" when X = 85 AND Y = 35 else
"111111111111" when X = 86 AND Y = 35 else
"111111111111" when X = 87 AND Y = 35 else
"111111111111" when X = 88 AND Y = 35 else
"111111111111" when X = 89 AND Y = 35 else
"111111111111" when X = 90 AND Y = 35 else
"111111111111" when X = 91 AND Y = 35 else
"111111111111" when X = 92 AND Y = 35 else
"111111111111" when X = 93 AND Y = 35 else
"111111111111" when X = 94 AND Y = 35 else
"111111111111" when X = 95 AND Y = 35 else
"111111111111" when X = 96 AND Y = 35 else
"111111111111" when X = 97 AND Y = 35 else
"111111111111" when X = 98 AND Y = 35 else
"111111111111" when X = 99 AND Y = 35 else
"111111111111" when X = 100 AND Y = 35 else
"111111111111" when X = 101 AND Y = 35 else
"111111111111" when X = 102 AND Y = 35 else
"111111111111" when X = 103 AND Y = 35 else
"111111111111" when X = 104 AND Y = 35 else
"111111111111" when X = 105 AND Y = 35 else
"111111111111" when X = 106 AND Y = 35 else
"111111111111" when X = 107 AND Y = 35 else
"111111111111" when X = 108 AND Y = 35 else
"111111111111" when X = 109 AND Y = 35 else
"111111111111" when X = 110 AND Y = 35 else
"111111111111" when X = 111 AND Y = 35 else
"111111111111" when X = 112 AND Y = 35 else
"111111111111" when X = 113 AND Y = 35 else
"111111111111" when X = 114 AND Y = 35 else
"111111111111" when X = 115 AND Y = 35 else
"111111111111" when X = 116 AND Y = 35 else
"111111111111" when X = 117 AND Y = 35 else
"111111111111" when X = 118 AND Y = 35 else
"111111111111" when X = 119 AND Y = 35 else
"111111111111" when X = 120 AND Y = 35 else
"111111111111" when X = 121 AND Y = 35 else
"111111111111" when X = 122 AND Y = 35 else
"111111111111" when X = 123 AND Y = 35 else
"111111111111" when X = 124 AND Y = 35 else
"111111111111" when X = 125 AND Y = 35 else
"111111111111" when X = 126 AND Y = 35 else
"111111111111" when X = 127 AND Y = 35 else
"111111111111" when X = 128 AND Y = 35 else
"111111111111" when X = 129 AND Y = 35 else
"111111111111" when X = 130 AND Y = 35 else
"111111111111" when X = 131 AND Y = 35 else
"111111111111" when X = 132 AND Y = 35 else
"111111111111" when X = 133 AND Y = 35 else
"111111111111" when X = 134 AND Y = 35 else
"111111111111" when X = 135 AND Y = 35 else
"111111111111" when X = 136 AND Y = 35 else
"111111111111" when X = 137 AND Y = 35 else
"111111111111" when X = 138 AND Y = 35 else
"111111111111" when X = 139 AND Y = 35 else
"111111111111" when X = 140 AND Y = 35 else
"111111111111" when X = 141 AND Y = 35 else
"111111111111" when X = 142 AND Y = 35 else
"111111111111" when X = 143 AND Y = 35 else
"111111111111" when X = 144 AND Y = 35 else
"111111111111" when X = 145 AND Y = 35 else
"111111111111" when X = 146 AND Y = 35 else
"111111111111" when X = 147 AND Y = 35 else
"111111111111" when X = 148 AND Y = 35 else
"111111111111" when X = 149 AND Y = 35 else
"111111111111" when X = 150 AND Y = 35 else
"111111111111" when X = 151 AND Y = 35 else
"111111111111" when X = 152 AND Y = 35 else
"111111111111" when X = 153 AND Y = 35 else
"111111111111" when X = 154 AND Y = 35 else
"111111111111" when X = 155 AND Y = 35 else
"111111111111" when X = 156 AND Y = 35 else
"111111111111" when X = 157 AND Y = 35 else
"111111111111" when X = 158 AND Y = 35 else
"111111111111" when X = 159 AND Y = 35 else
"111111111111" when X = 160 AND Y = 35 else
"111111111111" when X = 161 AND Y = 35 else
"111111111111" when X = 162 AND Y = 35 else
"111111111111" when X = 163 AND Y = 35 else
"111111111111" when X = 164 AND Y = 35 else
"111111111111" when X = 165 AND Y = 35 else
"111111111111" when X = 166 AND Y = 35 else
"111111111111" when X = 167 AND Y = 35 else
"111111111111" when X = 168 AND Y = 35 else
"111111111111" when X = 169 AND Y = 35 else
"111111111111" when X = 170 AND Y = 35 else
"111111111111" when X = 171 AND Y = 35 else
"111111111111" when X = 172 AND Y = 35 else
"111111111111" when X = 173 AND Y = 35 else
"111111111111" when X = 174 AND Y = 35 else
"111111111111" when X = 175 AND Y = 35 else
"111111111111" when X = 176 AND Y = 35 else
"111111111111" when X = 177 AND Y = 35 else
"111111111111" when X = 178 AND Y = 35 else
"111111111111" when X = 179 AND Y = 35 else
"111111111111" when X = 180 AND Y = 35 else
"111111111111" when X = 181 AND Y = 35 else
"111111111111" when X = 182 AND Y = 35 else
"111111111111" when X = 183 AND Y = 35 else
"111111111111" when X = 184 AND Y = 35 else
"111111111111" when X = 185 AND Y = 35 else
"111111111111" when X = 186 AND Y = 35 else
"111111111111" when X = 187 AND Y = 35 else
"111111111111" when X = 188 AND Y = 35 else
"111111111111" when X = 189 AND Y = 35 else
"111111111111" when X = 190 AND Y = 35 else
"111111111111" when X = 191 AND Y = 35 else
"111111111111" when X = 192 AND Y = 35 else
"111111111111" when X = 193 AND Y = 35 else
"111111111111" when X = 194 AND Y = 35 else
"111111111111" when X = 195 AND Y = 35 else
"111111111111" when X = 196 AND Y = 35 else
"111111111111" when X = 197 AND Y = 35 else
"111111111111" when X = 198 AND Y = 35 else
"111111111111" when X = 199 AND Y = 35 else
"000000000000" when X = 200 AND Y = 35 else
"000000000000" when X = 201 AND Y = 35 else
"000000000000" when X = 202 AND Y = 35 else
"000000000000" when X = 203 AND Y = 35 else
"000000000000" when X = 204 AND Y = 35 else
"000000000000" when X = 205 AND Y = 35 else
"000000000000" when X = 206 AND Y = 35 else
"000000000000" when X = 207 AND Y = 35 else
"000000000000" when X = 208 AND Y = 35 else
"000000000000" when X = 209 AND Y = 35 else
"000000000000" when X = 210 AND Y = 35 else
"000000000000" when X = 211 AND Y = 35 else
"000000000000" when X = 212 AND Y = 35 else
"000000000000" when X = 213 AND Y = 35 else
"000000000000" when X = 214 AND Y = 35 else
"111111111111" when X = 215 AND Y = 35 else
"111111111111" when X = 216 AND Y = 35 else
"111111111111" when X = 217 AND Y = 35 else
"111111111111" when X = 218 AND Y = 35 else
"111111111111" when X = 219 AND Y = 35 else
"111111111111" when X = 220 AND Y = 35 else
"111111111111" when X = 221 AND Y = 35 else
"111111111111" when X = 222 AND Y = 35 else
"111111111111" when X = 223 AND Y = 35 else
"111111111111" when X = 224 AND Y = 35 else
"111111111111" when X = 225 AND Y = 35 else
"111111111111" when X = 226 AND Y = 35 else
"111111111111" when X = 227 AND Y = 35 else
"111111111111" when X = 228 AND Y = 35 else
"111111111111" when X = 229 AND Y = 35 else
"111111111111" when X = 230 AND Y = 35 else
"111111111111" when X = 231 AND Y = 35 else
"111111111111" when X = 232 AND Y = 35 else
"111111111111" when X = 233 AND Y = 35 else
"111111111111" when X = 234 AND Y = 35 else
"111111111111" when X = 235 AND Y = 35 else
"111111111111" when X = 236 AND Y = 35 else
"111111111111" when X = 237 AND Y = 35 else
"111111111111" when X = 238 AND Y = 35 else
"111111111111" when X = 239 AND Y = 35 else
"111111111111" when X = 240 AND Y = 35 else
"111111111111" when X = 241 AND Y = 35 else
"111111111111" when X = 242 AND Y = 35 else
"111111111111" when X = 243 AND Y = 35 else
"111111111111" when X = 244 AND Y = 35 else
"111111111111" when X = 245 AND Y = 35 else
"111111111111" when X = 246 AND Y = 35 else
"111111111111" when X = 247 AND Y = 35 else
"111111111111" when X = 248 AND Y = 35 else
"111111111111" when X = 249 AND Y = 35 else
"111111111111" when X = 250 AND Y = 35 else
"111111111111" when X = 251 AND Y = 35 else
"111111111111" when X = 252 AND Y = 35 else
"111111111111" when X = 253 AND Y = 35 else
"111111111111" when X = 254 AND Y = 35 else
"111111111111" when X = 255 AND Y = 35 else
"111111111111" when X = 256 AND Y = 35 else
"111111111111" when X = 257 AND Y = 35 else
"111111111111" when X = 258 AND Y = 35 else
"111111111111" when X = 259 AND Y = 35 else
"110111011111" when X = 260 AND Y = 35 else
"110111011111" when X = 261 AND Y = 35 else
"110111011111" when X = 262 AND Y = 35 else
"110111011111" when X = 263 AND Y = 35 else
"110111011111" when X = 264 AND Y = 35 else
"110111011111" when X = 265 AND Y = 35 else
"110111011111" when X = 266 AND Y = 35 else
"110111011111" when X = 267 AND Y = 35 else
"110111011111" when X = 268 AND Y = 35 else
"110111011111" when X = 269 AND Y = 35 else
"110111011111" when X = 270 AND Y = 35 else
"110111011111" when X = 271 AND Y = 35 else
"110111011111" when X = 272 AND Y = 35 else
"110111011111" when X = 273 AND Y = 35 else
"110111011111" when X = 274 AND Y = 35 else
"110111011111" when X = 275 AND Y = 35 else
"110111011111" when X = 276 AND Y = 35 else
"110111011111" when X = 277 AND Y = 35 else
"110111011111" when X = 278 AND Y = 35 else
"110111011111" when X = 279 AND Y = 35 else
"000000000000" when X = 280 AND Y = 35 else
"000000000000" when X = 281 AND Y = 35 else
"000000000000" when X = 282 AND Y = 35 else
"000000000000" when X = 283 AND Y = 35 else
"000000000000" when X = 284 AND Y = 35 else
"000000000000" when X = 285 AND Y = 35 else
"000000000000" when X = 286 AND Y = 35 else
"000000000000" when X = 287 AND Y = 35 else
"000000000000" when X = 288 AND Y = 35 else
"000000000000" when X = 289 AND Y = 35 else
"000000000000" when X = 290 AND Y = 35 else
"000000000000" when X = 291 AND Y = 35 else
"000000000000" when X = 292 AND Y = 35 else
"000000000000" when X = 293 AND Y = 35 else
"000000000000" when X = 294 AND Y = 35 else
"000000000000" when X = 295 AND Y = 35 else
"000000000000" when X = 296 AND Y = 35 else
"000000000000" when X = 297 AND Y = 35 else
"000000000000" when X = 298 AND Y = 35 else
"000000000000" when X = 299 AND Y = 35 else
"000000000000" when X = 300 AND Y = 35 else
"000000000000" when X = 301 AND Y = 35 else
"000000000000" when X = 302 AND Y = 35 else
"000000000000" when X = 303 AND Y = 35 else
"000000000000" when X = 304 AND Y = 35 else
"000000000000" when X = 305 AND Y = 35 else
"000000000000" when X = 306 AND Y = 35 else
"000000000000" when X = 307 AND Y = 35 else
"000000000000" when X = 308 AND Y = 35 else
"000000000000" when X = 309 AND Y = 35 else
"000000000000" when X = 310 AND Y = 35 else
"000000000000" when X = 311 AND Y = 35 else
"000000000000" when X = 312 AND Y = 35 else
"000000000000" when X = 313 AND Y = 35 else
"000000000000" when X = 314 AND Y = 35 else
"000000000000" when X = 315 AND Y = 35 else
"000000000000" when X = 316 AND Y = 35 else
"000000000000" when X = 317 AND Y = 35 else
"000000000000" when X = 318 AND Y = 35 else
"000000000000" when X = 319 AND Y = 35 else
"000000000000" when X = 320 AND Y = 35 else
"000000000000" when X = 321 AND Y = 35 else
"000000000000" when X = 322 AND Y = 35 else
"000000000000" when X = 323 AND Y = 35 else
"000000000000" when X = 324 AND Y = 35 else
"000000000000" when X = 0 AND Y = 36 else
"000000000000" when X = 1 AND Y = 36 else
"000000000000" when X = 2 AND Y = 36 else
"000000000000" when X = 3 AND Y = 36 else
"000000000000" when X = 4 AND Y = 36 else
"000000000000" when X = 5 AND Y = 36 else
"000000000000" when X = 6 AND Y = 36 else
"000000000000" when X = 7 AND Y = 36 else
"000000000000" when X = 8 AND Y = 36 else
"000000000000" when X = 9 AND Y = 36 else
"000000000000" when X = 10 AND Y = 36 else
"000000000000" when X = 11 AND Y = 36 else
"000000000000" when X = 12 AND Y = 36 else
"000000000000" when X = 13 AND Y = 36 else
"000000000000" when X = 14 AND Y = 36 else
"000000000000" when X = 15 AND Y = 36 else
"000000000000" when X = 16 AND Y = 36 else
"000000000000" when X = 17 AND Y = 36 else
"000000000000" when X = 18 AND Y = 36 else
"000000000000" when X = 19 AND Y = 36 else
"000000000000" when X = 20 AND Y = 36 else
"000000000000" when X = 21 AND Y = 36 else
"000000000000" when X = 22 AND Y = 36 else
"000000000000" when X = 23 AND Y = 36 else
"000000000000" when X = 24 AND Y = 36 else
"000000000000" when X = 25 AND Y = 36 else
"000000000000" when X = 26 AND Y = 36 else
"000000000000" when X = 27 AND Y = 36 else
"000000000000" when X = 28 AND Y = 36 else
"000000000000" when X = 29 AND Y = 36 else
"000000000000" when X = 30 AND Y = 36 else
"000000000000" when X = 31 AND Y = 36 else
"000000000000" when X = 32 AND Y = 36 else
"000000000000" when X = 33 AND Y = 36 else
"000000000000" when X = 34 AND Y = 36 else
"000000000000" when X = 35 AND Y = 36 else
"000000000000" when X = 36 AND Y = 36 else
"000000000000" when X = 37 AND Y = 36 else
"000000000000" when X = 38 AND Y = 36 else
"000000000000" when X = 39 AND Y = 36 else
"100010011101" when X = 40 AND Y = 36 else
"100010011101" when X = 41 AND Y = 36 else
"100010011101" when X = 42 AND Y = 36 else
"100010011101" when X = 43 AND Y = 36 else
"100010011101" when X = 44 AND Y = 36 else
"100010011101" when X = 45 AND Y = 36 else
"100010011101" when X = 46 AND Y = 36 else
"100010011101" when X = 47 AND Y = 36 else
"100010011101" when X = 48 AND Y = 36 else
"100010011101" when X = 49 AND Y = 36 else
"110111011111" when X = 50 AND Y = 36 else
"110111011111" when X = 51 AND Y = 36 else
"110111011111" when X = 52 AND Y = 36 else
"110111011111" when X = 53 AND Y = 36 else
"110111011111" when X = 54 AND Y = 36 else
"110111011111" when X = 55 AND Y = 36 else
"110111011111" when X = 56 AND Y = 36 else
"110111011111" when X = 57 AND Y = 36 else
"110111011111" when X = 58 AND Y = 36 else
"110111011111" when X = 59 AND Y = 36 else
"111111111111" when X = 60 AND Y = 36 else
"111111111111" when X = 61 AND Y = 36 else
"111111111111" when X = 62 AND Y = 36 else
"111111111111" when X = 63 AND Y = 36 else
"111111111111" when X = 64 AND Y = 36 else
"111111111111" when X = 65 AND Y = 36 else
"111111111111" when X = 66 AND Y = 36 else
"111111111111" when X = 67 AND Y = 36 else
"111111111111" when X = 68 AND Y = 36 else
"111111111111" when X = 69 AND Y = 36 else
"111111111111" when X = 70 AND Y = 36 else
"111111111111" when X = 71 AND Y = 36 else
"111111111111" when X = 72 AND Y = 36 else
"111111111111" when X = 73 AND Y = 36 else
"111111111111" when X = 74 AND Y = 36 else
"111111111111" when X = 75 AND Y = 36 else
"111111111111" when X = 76 AND Y = 36 else
"111111111111" when X = 77 AND Y = 36 else
"111111111111" when X = 78 AND Y = 36 else
"111111111111" when X = 79 AND Y = 36 else
"111111111111" when X = 80 AND Y = 36 else
"111111111111" when X = 81 AND Y = 36 else
"111111111111" when X = 82 AND Y = 36 else
"111111111111" when X = 83 AND Y = 36 else
"111111111111" when X = 84 AND Y = 36 else
"111111111111" when X = 85 AND Y = 36 else
"111111111111" when X = 86 AND Y = 36 else
"111111111111" when X = 87 AND Y = 36 else
"111111111111" when X = 88 AND Y = 36 else
"111111111111" when X = 89 AND Y = 36 else
"111111111111" when X = 90 AND Y = 36 else
"111111111111" when X = 91 AND Y = 36 else
"111111111111" when X = 92 AND Y = 36 else
"111111111111" when X = 93 AND Y = 36 else
"111111111111" when X = 94 AND Y = 36 else
"111111111111" when X = 95 AND Y = 36 else
"111111111111" when X = 96 AND Y = 36 else
"111111111111" when X = 97 AND Y = 36 else
"111111111111" when X = 98 AND Y = 36 else
"111111111111" when X = 99 AND Y = 36 else
"111111111111" when X = 100 AND Y = 36 else
"111111111111" when X = 101 AND Y = 36 else
"111111111111" when X = 102 AND Y = 36 else
"111111111111" when X = 103 AND Y = 36 else
"111111111111" when X = 104 AND Y = 36 else
"111111111111" when X = 105 AND Y = 36 else
"111111111111" when X = 106 AND Y = 36 else
"111111111111" when X = 107 AND Y = 36 else
"111111111111" when X = 108 AND Y = 36 else
"111111111111" when X = 109 AND Y = 36 else
"111111111111" when X = 110 AND Y = 36 else
"111111111111" when X = 111 AND Y = 36 else
"111111111111" when X = 112 AND Y = 36 else
"111111111111" when X = 113 AND Y = 36 else
"111111111111" when X = 114 AND Y = 36 else
"111111111111" when X = 115 AND Y = 36 else
"111111111111" when X = 116 AND Y = 36 else
"111111111111" when X = 117 AND Y = 36 else
"111111111111" when X = 118 AND Y = 36 else
"111111111111" when X = 119 AND Y = 36 else
"111111111111" when X = 120 AND Y = 36 else
"111111111111" when X = 121 AND Y = 36 else
"111111111111" when X = 122 AND Y = 36 else
"111111111111" when X = 123 AND Y = 36 else
"111111111111" when X = 124 AND Y = 36 else
"111111111111" when X = 125 AND Y = 36 else
"111111111111" when X = 126 AND Y = 36 else
"111111111111" when X = 127 AND Y = 36 else
"111111111111" when X = 128 AND Y = 36 else
"111111111111" when X = 129 AND Y = 36 else
"111111111111" when X = 130 AND Y = 36 else
"111111111111" when X = 131 AND Y = 36 else
"111111111111" when X = 132 AND Y = 36 else
"111111111111" when X = 133 AND Y = 36 else
"111111111111" when X = 134 AND Y = 36 else
"111111111111" when X = 135 AND Y = 36 else
"111111111111" when X = 136 AND Y = 36 else
"111111111111" when X = 137 AND Y = 36 else
"111111111111" when X = 138 AND Y = 36 else
"111111111111" when X = 139 AND Y = 36 else
"111111111111" when X = 140 AND Y = 36 else
"111111111111" when X = 141 AND Y = 36 else
"111111111111" when X = 142 AND Y = 36 else
"111111111111" when X = 143 AND Y = 36 else
"111111111111" when X = 144 AND Y = 36 else
"111111111111" when X = 145 AND Y = 36 else
"111111111111" when X = 146 AND Y = 36 else
"111111111111" when X = 147 AND Y = 36 else
"111111111111" when X = 148 AND Y = 36 else
"111111111111" when X = 149 AND Y = 36 else
"111111111111" when X = 150 AND Y = 36 else
"111111111111" when X = 151 AND Y = 36 else
"111111111111" when X = 152 AND Y = 36 else
"111111111111" when X = 153 AND Y = 36 else
"111111111111" when X = 154 AND Y = 36 else
"111111111111" when X = 155 AND Y = 36 else
"111111111111" when X = 156 AND Y = 36 else
"111111111111" when X = 157 AND Y = 36 else
"111111111111" when X = 158 AND Y = 36 else
"111111111111" when X = 159 AND Y = 36 else
"111111111111" when X = 160 AND Y = 36 else
"111111111111" when X = 161 AND Y = 36 else
"111111111111" when X = 162 AND Y = 36 else
"111111111111" when X = 163 AND Y = 36 else
"111111111111" when X = 164 AND Y = 36 else
"111111111111" when X = 165 AND Y = 36 else
"111111111111" when X = 166 AND Y = 36 else
"111111111111" when X = 167 AND Y = 36 else
"111111111111" when X = 168 AND Y = 36 else
"111111111111" when X = 169 AND Y = 36 else
"111111111111" when X = 170 AND Y = 36 else
"111111111111" when X = 171 AND Y = 36 else
"111111111111" when X = 172 AND Y = 36 else
"111111111111" when X = 173 AND Y = 36 else
"111111111111" when X = 174 AND Y = 36 else
"111111111111" when X = 175 AND Y = 36 else
"111111111111" when X = 176 AND Y = 36 else
"111111111111" when X = 177 AND Y = 36 else
"111111111111" when X = 178 AND Y = 36 else
"111111111111" when X = 179 AND Y = 36 else
"111111111111" when X = 180 AND Y = 36 else
"111111111111" when X = 181 AND Y = 36 else
"111111111111" when X = 182 AND Y = 36 else
"111111111111" when X = 183 AND Y = 36 else
"111111111111" when X = 184 AND Y = 36 else
"111111111111" when X = 185 AND Y = 36 else
"111111111111" when X = 186 AND Y = 36 else
"111111111111" when X = 187 AND Y = 36 else
"111111111111" when X = 188 AND Y = 36 else
"111111111111" when X = 189 AND Y = 36 else
"111111111111" when X = 190 AND Y = 36 else
"111111111111" when X = 191 AND Y = 36 else
"111111111111" when X = 192 AND Y = 36 else
"111111111111" when X = 193 AND Y = 36 else
"111111111111" when X = 194 AND Y = 36 else
"111111111111" when X = 195 AND Y = 36 else
"111111111111" when X = 196 AND Y = 36 else
"111111111111" when X = 197 AND Y = 36 else
"111111111111" when X = 198 AND Y = 36 else
"111111111111" when X = 199 AND Y = 36 else
"000000000000" when X = 200 AND Y = 36 else
"000000000000" when X = 201 AND Y = 36 else
"000000000000" when X = 202 AND Y = 36 else
"000000000000" when X = 203 AND Y = 36 else
"000000000000" when X = 204 AND Y = 36 else
"000000000000" when X = 205 AND Y = 36 else
"000000000000" when X = 206 AND Y = 36 else
"000000000000" when X = 207 AND Y = 36 else
"000000000000" when X = 208 AND Y = 36 else
"000000000000" when X = 209 AND Y = 36 else
"000000000000" when X = 210 AND Y = 36 else
"000000000000" when X = 211 AND Y = 36 else
"000000000000" when X = 212 AND Y = 36 else
"000000000000" when X = 213 AND Y = 36 else
"000000000000" when X = 214 AND Y = 36 else
"111111111111" when X = 215 AND Y = 36 else
"111111111111" when X = 216 AND Y = 36 else
"111111111111" when X = 217 AND Y = 36 else
"111111111111" when X = 218 AND Y = 36 else
"111111111111" when X = 219 AND Y = 36 else
"111111111111" when X = 220 AND Y = 36 else
"111111111111" when X = 221 AND Y = 36 else
"111111111111" when X = 222 AND Y = 36 else
"111111111111" when X = 223 AND Y = 36 else
"111111111111" when X = 224 AND Y = 36 else
"111111111111" when X = 225 AND Y = 36 else
"111111111111" when X = 226 AND Y = 36 else
"111111111111" when X = 227 AND Y = 36 else
"111111111111" when X = 228 AND Y = 36 else
"111111111111" when X = 229 AND Y = 36 else
"111111111111" when X = 230 AND Y = 36 else
"111111111111" when X = 231 AND Y = 36 else
"111111111111" when X = 232 AND Y = 36 else
"111111111111" when X = 233 AND Y = 36 else
"111111111111" when X = 234 AND Y = 36 else
"111111111111" when X = 235 AND Y = 36 else
"111111111111" when X = 236 AND Y = 36 else
"111111111111" when X = 237 AND Y = 36 else
"111111111111" when X = 238 AND Y = 36 else
"111111111111" when X = 239 AND Y = 36 else
"111111111111" when X = 240 AND Y = 36 else
"111111111111" when X = 241 AND Y = 36 else
"111111111111" when X = 242 AND Y = 36 else
"111111111111" when X = 243 AND Y = 36 else
"111111111111" when X = 244 AND Y = 36 else
"111111111111" when X = 245 AND Y = 36 else
"111111111111" when X = 246 AND Y = 36 else
"111111111111" when X = 247 AND Y = 36 else
"111111111111" when X = 248 AND Y = 36 else
"111111111111" when X = 249 AND Y = 36 else
"111111111111" when X = 250 AND Y = 36 else
"111111111111" when X = 251 AND Y = 36 else
"111111111111" when X = 252 AND Y = 36 else
"111111111111" when X = 253 AND Y = 36 else
"111111111111" when X = 254 AND Y = 36 else
"111111111111" when X = 255 AND Y = 36 else
"111111111111" when X = 256 AND Y = 36 else
"111111111111" when X = 257 AND Y = 36 else
"111111111111" when X = 258 AND Y = 36 else
"111111111111" when X = 259 AND Y = 36 else
"110111011111" when X = 260 AND Y = 36 else
"110111011111" when X = 261 AND Y = 36 else
"110111011111" when X = 262 AND Y = 36 else
"110111011111" when X = 263 AND Y = 36 else
"110111011111" when X = 264 AND Y = 36 else
"110111011111" when X = 265 AND Y = 36 else
"110111011111" when X = 266 AND Y = 36 else
"110111011111" when X = 267 AND Y = 36 else
"110111011111" when X = 268 AND Y = 36 else
"110111011111" when X = 269 AND Y = 36 else
"110111011111" when X = 270 AND Y = 36 else
"110111011111" when X = 271 AND Y = 36 else
"110111011111" when X = 272 AND Y = 36 else
"110111011111" when X = 273 AND Y = 36 else
"110111011111" when X = 274 AND Y = 36 else
"110111011111" when X = 275 AND Y = 36 else
"110111011111" when X = 276 AND Y = 36 else
"110111011111" when X = 277 AND Y = 36 else
"110111011111" when X = 278 AND Y = 36 else
"110111011111" when X = 279 AND Y = 36 else
"000000000000" when X = 280 AND Y = 36 else
"000000000000" when X = 281 AND Y = 36 else
"000000000000" when X = 282 AND Y = 36 else
"000000000000" when X = 283 AND Y = 36 else
"000000000000" when X = 284 AND Y = 36 else
"000000000000" when X = 285 AND Y = 36 else
"000000000000" when X = 286 AND Y = 36 else
"000000000000" when X = 287 AND Y = 36 else
"000000000000" when X = 288 AND Y = 36 else
"000000000000" when X = 289 AND Y = 36 else
"000000000000" when X = 290 AND Y = 36 else
"000000000000" when X = 291 AND Y = 36 else
"000000000000" when X = 292 AND Y = 36 else
"000000000000" when X = 293 AND Y = 36 else
"000000000000" when X = 294 AND Y = 36 else
"000000000000" when X = 295 AND Y = 36 else
"000000000000" when X = 296 AND Y = 36 else
"000000000000" when X = 297 AND Y = 36 else
"000000000000" when X = 298 AND Y = 36 else
"000000000000" when X = 299 AND Y = 36 else
"000000000000" when X = 300 AND Y = 36 else
"000000000000" when X = 301 AND Y = 36 else
"000000000000" when X = 302 AND Y = 36 else
"000000000000" when X = 303 AND Y = 36 else
"000000000000" when X = 304 AND Y = 36 else
"000000000000" when X = 305 AND Y = 36 else
"000000000000" when X = 306 AND Y = 36 else
"000000000000" when X = 307 AND Y = 36 else
"000000000000" when X = 308 AND Y = 36 else
"000000000000" when X = 309 AND Y = 36 else
"000000000000" when X = 310 AND Y = 36 else
"000000000000" when X = 311 AND Y = 36 else
"000000000000" when X = 312 AND Y = 36 else
"000000000000" when X = 313 AND Y = 36 else
"000000000000" when X = 314 AND Y = 36 else
"000000000000" when X = 315 AND Y = 36 else
"000000000000" when X = 316 AND Y = 36 else
"000000000000" when X = 317 AND Y = 36 else
"000000000000" when X = 318 AND Y = 36 else
"000000000000" when X = 319 AND Y = 36 else
"000000000000" when X = 320 AND Y = 36 else
"000000000000" when X = 321 AND Y = 36 else
"000000000000" when X = 322 AND Y = 36 else
"000000000000" when X = 323 AND Y = 36 else
"000000000000" when X = 324 AND Y = 36 else
"000000000000" when X = 0 AND Y = 37 else
"000000000000" when X = 1 AND Y = 37 else
"000000000000" when X = 2 AND Y = 37 else
"000000000000" when X = 3 AND Y = 37 else
"000000000000" when X = 4 AND Y = 37 else
"000000000000" when X = 5 AND Y = 37 else
"000000000000" when X = 6 AND Y = 37 else
"000000000000" when X = 7 AND Y = 37 else
"000000000000" when X = 8 AND Y = 37 else
"000000000000" when X = 9 AND Y = 37 else
"000000000000" when X = 10 AND Y = 37 else
"000000000000" when X = 11 AND Y = 37 else
"000000000000" when X = 12 AND Y = 37 else
"000000000000" when X = 13 AND Y = 37 else
"000000000000" when X = 14 AND Y = 37 else
"000000000000" when X = 15 AND Y = 37 else
"000000000000" when X = 16 AND Y = 37 else
"000000000000" when X = 17 AND Y = 37 else
"000000000000" when X = 18 AND Y = 37 else
"000000000000" when X = 19 AND Y = 37 else
"000000000000" when X = 20 AND Y = 37 else
"000000000000" when X = 21 AND Y = 37 else
"000000000000" when X = 22 AND Y = 37 else
"000000000000" when X = 23 AND Y = 37 else
"000000000000" when X = 24 AND Y = 37 else
"000000000000" when X = 25 AND Y = 37 else
"000000000000" when X = 26 AND Y = 37 else
"000000000000" when X = 27 AND Y = 37 else
"000000000000" when X = 28 AND Y = 37 else
"000000000000" when X = 29 AND Y = 37 else
"000000000000" when X = 30 AND Y = 37 else
"000000000000" when X = 31 AND Y = 37 else
"000000000000" when X = 32 AND Y = 37 else
"000000000000" when X = 33 AND Y = 37 else
"000000000000" when X = 34 AND Y = 37 else
"000000000000" when X = 35 AND Y = 37 else
"000000000000" when X = 36 AND Y = 37 else
"000000000000" when X = 37 AND Y = 37 else
"000000000000" when X = 38 AND Y = 37 else
"000000000000" when X = 39 AND Y = 37 else
"100010011101" when X = 40 AND Y = 37 else
"100010011101" when X = 41 AND Y = 37 else
"100010011101" when X = 42 AND Y = 37 else
"100010011101" when X = 43 AND Y = 37 else
"100010011101" when X = 44 AND Y = 37 else
"100010011101" when X = 45 AND Y = 37 else
"100010011101" when X = 46 AND Y = 37 else
"100010011101" when X = 47 AND Y = 37 else
"100010011101" when X = 48 AND Y = 37 else
"100010011101" when X = 49 AND Y = 37 else
"110111011111" when X = 50 AND Y = 37 else
"110111011111" when X = 51 AND Y = 37 else
"110111011111" when X = 52 AND Y = 37 else
"110111011111" when X = 53 AND Y = 37 else
"110111011111" when X = 54 AND Y = 37 else
"110111011111" when X = 55 AND Y = 37 else
"110111011111" when X = 56 AND Y = 37 else
"110111011111" when X = 57 AND Y = 37 else
"110111011111" when X = 58 AND Y = 37 else
"110111011111" when X = 59 AND Y = 37 else
"111111111111" when X = 60 AND Y = 37 else
"111111111111" when X = 61 AND Y = 37 else
"111111111111" when X = 62 AND Y = 37 else
"111111111111" when X = 63 AND Y = 37 else
"111111111111" when X = 64 AND Y = 37 else
"111111111111" when X = 65 AND Y = 37 else
"111111111111" when X = 66 AND Y = 37 else
"111111111111" when X = 67 AND Y = 37 else
"111111111111" when X = 68 AND Y = 37 else
"111111111111" when X = 69 AND Y = 37 else
"111111111111" when X = 70 AND Y = 37 else
"111111111111" when X = 71 AND Y = 37 else
"111111111111" when X = 72 AND Y = 37 else
"111111111111" when X = 73 AND Y = 37 else
"111111111111" when X = 74 AND Y = 37 else
"111111111111" when X = 75 AND Y = 37 else
"111111111111" when X = 76 AND Y = 37 else
"111111111111" when X = 77 AND Y = 37 else
"111111111111" when X = 78 AND Y = 37 else
"111111111111" when X = 79 AND Y = 37 else
"111111111111" when X = 80 AND Y = 37 else
"111111111111" when X = 81 AND Y = 37 else
"111111111111" when X = 82 AND Y = 37 else
"111111111111" when X = 83 AND Y = 37 else
"111111111111" when X = 84 AND Y = 37 else
"111111111111" when X = 85 AND Y = 37 else
"111111111111" when X = 86 AND Y = 37 else
"111111111111" when X = 87 AND Y = 37 else
"111111111111" when X = 88 AND Y = 37 else
"111111111111" when X = 89 AND Y = 37 else
"111111111111" when X = 90 AND Y = 37 else
"111111111111" when X = 91 AND Y = 37 else
"111111111111" when X = 92 AND Y = 37 else
"111111111111" when X = 93 AND Y = 37 else
"111111111111" when X = 94 AND Y = 37 else
"111111111111" when X = 95 AND Y = 37 else
"111111111111" when X = 96 AND Y = 37 else
"111111111111" when X = 97 AND Y = 37 else
"111111111111" when X = 98 AND Y = 37 else
"111111111111" when X = 99 AND Y = 37 else
"111111111111" when X = 100 AND Y = 37 else
"111111111111" when X = 101 AND Y = 37 else
"111111111111" when X = 102 AND Y = 37 else
"111111111111" when X = 103 AND Y = 37 else
"111111111111" when X = 104 AND Y = 37 else
"111111111111" when X = 105 AND Y = 37 else
"111111111111" when X = 106 AND Y = 37 else
"111111111111" when X = 107 AND Y = 37 else
"111111111111" when X = 108 AND Y = 37 else
"111111111111" when X = 109 AND Y = 37 else
"111111111111" when X = 110 AND Y = 37 else
"111111111111" when X = 111 AND Y = 37 else
"111111111111" when X = 112 AND Y = 37 else
"111111111111" when X = 113 AND Y = 37 else
"111111111111" when X = 114 AND Y = 37 else
"111111111111" when X = 115 AND Y = 37 else
"111111111111" when X = 116 AND Y = 37 else
"111111111111" when X = 117 AND Y = 37 else
"111111111111" when X = 118 AND Y = 37 else
"111111111111" when X = 119 AND Y = 37 else
"111111111111" when X = 120 AND Y = 37 else
"111111111111" when X = 121 AND Y = 37 else
"111111111111" when X = 122 AND Y = 37 else
"111111111111" when X = 123 AND Y = 37 else
"111111111111" when X = 124 AND Y = 37 else
"111111111111" when X = 125 AND Y = 37 else
"111111111111" when X = 126 AND Y = 37 else
"111111111111" when X = 127 AND Y = 37 else
"111111111111" when X = 128 AND Y = 37 else
"111111111111" when X = 129 AND Y = 37 else
"111111111111" when X = 130 AND Y = 37 else
"111111111111" when X = 131 AND Y = 37 else
"111111111111" when X = 132 AND Y = 37 else
"111111111111" when X = 133 AND Y = 37 else
"111111111111" when X = 134 AND Y = 37 else
"111111111111" when X = 135 AND Y = 37 else
"111111111111" when X = 136 AND Y = 37 else
"111111111111" when X = 137 AND Y = 37 else
"111111111111" when X = 138 AND Y = 37 else
"111111111111" when X = 139 AND Y = 37 else
"111111111111" when X = 140 AND Y = 37 else
"111111111111" when X = 141 AND Y = 37 else
"111111111111" when X = 142 AND Y = 37 else
"111111111111" when X = 143 AND Y = 37 else
"111111111111" when X = 144 AND Y = 37 else
"111111111111" when X = 145 AND Y = 37 else
"111111111111" when X = 146 AND Y = 37 else
"111111111111" when X = 147 AND Y = 37 else
"111111111111" when X = 148 AND Y = 37 else
"111111111111" when X = 149 AND Y = 37 else
"111111111111" when X = 150 AND Y = 37 else
"111111111111" when X = 151 AND Y = 37 else
"111111111111" when X = 152 AND Y = 37 else
"111111111111" when X = 153 AND Y = 37 else
"111111111111" when X = 154 AND Y = 37 else
"111111111111" when X = 155 AND Y = 37 else
"111111111111" when X = 156 AND Y = 37 else
"111111111111" when X = 157 AND Y = 37 else
"111111111111" when X = 158 AND Y = 37 else
"111111111111" when X = 159 AND Y = 37 else
"111111111111" when X = 160 AND Y = 37 else
"111111111111" when X = 161 AND Y = 37 else
"111111111111" when X = 162 AND Y = 37 else
"111111111111" when X = 163 AND Y = 37 else
"111111111111" when X = 164 AND Y = 37 else
"111111111111" when X = 165 AND Y = 37 else
"111111111111" when X = 166 AND Y = 37 else
"111111111111" when X = 167 AND Y = 37 else
"111111111111" when X = 168 AND Y = 37 else
"111111111111" when X = 169 AND Y = 37 else
"111111111111" when X = 170 AND Y = 37 else
"111111111111" when X = 171 AND Y = 37 else
"111111111111" when X = 172 AND Y = 37 else
"111111111111" when X = 173 AND Y = 37 else
"111111111111" when X = 174 AND Y = 37 else
"111111111111" when X = 175 AND Y = 37 else
"111111111111" when X = 176 AND Y = 37 else
"111111111111" when X = 177 AND Y = 37 else
"111111111111" when X = 178 AND Y = 37 else
"111111111111" when X = 179 AND Y = 37 else
"111111111111" when X = 180 AND Y = 37 else
"111111111111" when X = 181 AND Y = 37 else
"111111111111" when X = 182 AND Y = 37 else
"111111111111" when X = 183 AND Y = 37 else
"111111111111" when X = 184 AND Y = 37 else
"111111111111" when X = 185 AND Y = 37 else
"111111111111" when X = 186 AND Y = 37 else
"111111111111" when X = 187 AND Y = 37 else
"111111111111" when X = 188 AND Y = 37 else
"111111111111" when X = 189 AND Y = 37 else
"111111111111" when X = 190 AND Y = 37 else
"111111111111" when X = 191 AND Y = 37 else
"111111111111" when X = 192 AND Y = 37 else
"111111111111" when X = 193 AND Y = 37 else
"111111111111" when X = 194 AND Y = 37 else
"111111111111" when X = 195 AND Y = 37 else
"111111111111" when X = 196 AND Y = 37 else
"111111111111" when X = 197 AND Y = 37 else
"111111111111" when X = 198 AND Y = 37 else
"111111111111" when X = 199 AND Y = 37 else
"000000000000" when X = 200 AND Y = 37 else
"000000000000" when X = 201 AND Y = 37 else
"000000000000" when X = 202 AND Y = 37 else
"000000000000" when X = 203 AND Y = 37 else
"000000000000" when X = 204 AND Y = 37 else
"000000000000" when X = 205 AND Y = 37 else
"000000000000" when X = 206 AND Y = 37 else
"000000000000" when X = 207 AND Y = 37 else
"000000000000" when X = 208 AND Y = 37 else
"000000000000" when X = 209 AND Y = 37 else
"000000000000" when X = 210 AND Y = 37 else
"000000000000" when X = 211 AND Y = 37 else
"000000000000" when X = 212 AND Y = 37 else
"000000000000" when X = 213 AND Y = 37 else
"000000000000" when X = 214 AND Y = 37 else
"111111111111" when X = 215 AND Y = 37 else
"111111111111" when X = 216 AND Y = 37 else
"111111111111" when X = 217 AND Y = 37 else
"111111111111" when X = 218 AND Y = 37 else
"111111111111" when X = 219 AND Y = 37 else
"111111111111" when X = 220 AND Y = 37 else
"111111111111" when X = 221 AND Y = 37 else
"111111111111" when X = 222 AND Y = 37 else
"111111111111" when X = 223 AND Y = 37 else
"111111111111" when X = 224 AND Y = 37 else
"111111111111" when X = 225 AND Y = 37 else
"111111111111" when X = 226 AND Y = 37 else
"111111111111" when X = 227 AND Y = 37 else
"111111111111" when X = 228 AND Y = 37 else
"111111111111" when X = 229 AND Y = 37 else
"111111111111" when X = 230 AND Y = 37 else
"111111111111" when X = 231 AND Y = 37 else
"111111111111" when X = 232 AND Y = 37 else
"111111111111" when X = 233 AND Y = 37 else
"111111111111" when X = 234 AND Y = 37 else
"111111111111" when X = 235 AND Y = 37 else
"111111111111" when X = 236 AND Y = 37 else
"111111111111" when X = 237 AND Y = 37 else
"111111111111" when X = 238 AND Y = 37 else
"111111111111" when X = 239 AND Y = 37 else
"111111111111" when X = 240 AND Y = 37 else
"111111111111" when X = 241 AND Y = 37 else
"111111111111" when X = 242 AND Y = 37 else
"111111111111" when X = 243 AND Y = 37 else
"111111111111" when X = 244 AND Y = 37 else
"111111111111" when X = 245 AND Y = 37 else
"111111111111" when X = 246 AND Y = 37 else
"111111111111" when X = 247 AND Y = 37 else
"111111111111" when X = 248 AND Y = 37 else
"111111111111" when X = 249 AND Y = 37 else
"111111111111" when X = 250 AND Y = 37 else
"111111111111" when X = 251 AND Y = 37 else
"111111111111" when X = 252 AND Y = 37 else
"111111111111" when X = 253 AND Y = 37 else
"111111111111" when X = 254 AND Y = 37 else
"111111111111" when X = 255 AND Y = 37 else
"111111111111" when X = 256 AND Y = 37 else
"111111111111" when X = 257 AND Y = 37 else
"111111111111" when X = 258 AND Y = 37 else
"111111111111" when X = 259 AND Y = 37 else
"110111011111" when X = 260 AND Y = 37 else
"110111011111" when X = 261 AND Y = 37 else
"110111011111" when X = 262 AND Y = 37 else
"110111011111" when X = 263 AND Y = 37 else
"110111011111" when X = 264 AND Y = 37 else
"110111011111" when X = 265 AND Y = 37 else
"110111011111" when X = 266 AND Y = 37 else
"110111011111" when X = 267 AND Y = 37 else
"110111011111" when X = 268 AND Y = 37 else
"110111011111" when X = 269 AND Y = 37 else
"110111011111" when X = 270 AND Y = 37 else
"110111011111" when X = 271 AND Y = 37 else
"110111011111" when X = 272 AND Y = 37 else
"110111011111" when X = 273 AND Y = 37 else
"110111011111" when X = 274 AND Y = 37 else
"110111011111" when X = 275 AND Y = 37 else
"110111011111" when X = 276 AND Y = 37 else
"110111011111" when X = 277 AND Y = 37 else
"110111011111" when X = 278 AND Y = 37 else
"110111011111" when X = 279 AND Y = 37 else
"000000000000" when X = 280 AND Y = 37 else
"000000000000" when X = 281 AND Y = 37 else
"000000000000" when X = 282 AND Y = 37 else
"000000000000" when X = 283 AND Y = 37 else
"000000000000" when X = 284 AND Y = 37 else
"000000000000" when X = 285 AND Y = 37 else
"000000000000" when X = 286 AND Y = 37 else
"000000000000" when X = 287 AND Y = 37 else
"000000000000" when X = 288 AND Y = 37 else
"000000000000" when X = 289 AND Y = 37 else
"000000000000" when X = 290 AND Y = 37 else
"000000000000" when X = 291 AND Y = 37 else
"000000000000" when X = 292 AND Y = 37 else
"000000000000" when X = 293 AND Y = 37 else
"000000000000" when X = 294 AND Y = 37 else
"000000000000" when X = 295 AND Y = 37 else
"000000000000" when X = 296 AND Y = 37 else
"000000000000" when X = 297 AND Y = 37 else
"000000000000" when X = 298 AND Y = 37 else
"000000000000" when X = 299 AND Y = 37 else
"000000000000" when X = 300 AND Y = 37 else
"000000000000" when X = 301 AND Y = 37 else
"000000000000" when X = 302 AND Y = 37 else
"000000000000" when X = 303 AND Y = 37 else
"000000000000" when X = 304 AND Y = 37 else
"000000000000" when X = 305 AND Y = 37 else
"000000000000" when X = 306 AND Y = 37 else
"000000000000" when X = 307 AND Y = 37 else
"000000000000" when X = 308 AND Y = 37 else
"000000000000" when X = 309 AND Y = 37 else
"000000000000" when X = 310 AND Y = 37 else
"000000000000" when X = 311 AND Y = 37 else
"000000000000" when X = 312 AND Y = 37 else
"000000000000" when X = 313 AND Y = 37 else
"000000000000" when X = 314 AND Y = 37 else
"000000000000" when X = 315 AND Y = 37 else
"000000000000" when X = 316 AND Y = 37 else
"000000000000" when X = 317 AND Y = 37 else
"000000000000" when X = 318 AND Y = 37 else
"000000000000" when X = 319 AND Y = 37 else
"000000000000" when X = 320 AND Y = 37 else
"000000000000" when X = 321 AND Y = 37 else
"000000000000" when X = 322 AND Y = 37 else
"000000000000" when X = 323 AND Y = 37 else
"000000000000" when X = 324 AND Y = 37 else
"000000000000" when X = 0 AND Y = 38 else
"000000000000" when X = 1 AND Y = 38 else
"000000000000" when X = 2 AND Y = 38 else
"000000000000" when X = 3 AND Y = 38 else
"000000000000" when X = 4 AND Y = 38 else
"000000000000" when X = 5 AND Y = 38 else
"000000000000" when X = 6 AND Y = 38 else
"000000000000" when X = 7 AND Y = 38 else
"000000000000" when X = 8 AND Y = 38 else
"000000000000" when X = 9 AND Y = 38 else
"000000000000" when X = 10 AND Y = 38 else
"000000000000" when X = 11 AND Y = 38 else
"000000000000" when X = 12 AND Y = 38 else
"000000000000" when X = 13 AND Y = 38 else
"000000000000" when X = 14 AND Y = 38 else
"000000000000" when X = 15 AND Y = 38 else
"000000000000" when X = 16 AND Y = 38 else
"000000000000" when X = 17 AND Y = 38 else
"000000000000" when X = 18 AND Y = 38 else
"000000000000" when X = 19 AND Y = 38 else
"000000000000" when X = 20 AND Y = 38 else
"000000000000" when X = 21 AND Y = 38 else
"000000000000" when X = 22 AND Y = 38 else
"000000000000" when X = 23 AND Y = 38 else
"000000000000" when X = 24 AND Y = 38 else
"000000000000" when X = 25 AND Y = 38 else
"000000000000" when X = 26 AND Y = 38 else
"000000000000" when X = 27 AND Y = 38 else
"000000000000" when X = 28 AND Y = 38 else
"000000000000" when X = 29 AND Y = 38 else
"000000000000" when X = 30 AND Y = 38 else
"000000000000" when X = 31 AND Y = 38 else
"000000000000" when X = 32 AND Y = 38 else
"000000000000" when X = 33 AND Y = 38 else
"000000000000" when X = 34 AND Y = 38 else
"000000000000" when X = 35 AND Y = 38 else
"000000000000" when X = 36 AND Y = 38 else
"000000000000" when X = 37 AND Y = 38 else
"000000000000" when X = 38 AND Y = 38 else
"000000000000" when X = 39 AND Y = 38 else
"100010011101" when X = 40 AND Y = 38 else
"100010011101" when X = 41 AND Y = 38 else
"100010011101" when X = 42 AND Y = 38 else
"100010011101" when X = 43 AND Y = 38 else
"100010011101" when X = 44 AND Y = 38 else
"100010011101" when X = 45 AND Y = 38 else
"100010011101" when X = 46 AND Y = 38 else
"100010011101" when X = 47 AND Y = 38 else
"100010011101" when X = 48 AND Y = 38 else
"100010011101" when X = 49 AND Y = 38 else
"110111011111" when X = 50 AND Y = 38 else
"110111011111" when X = 51 AND Y = 38 else
"110111011111" when X = 52 AND Y = 38 else
"110111011111" when X = 53 AND Y = 38 else
"110111011111" when X = 54 AND Y = 38 else
"110111011111" when X = 55 AND Y = 38 else
"110111011111" when X = 56 AND Y = 38 else
"110111011111" when X = 57 AND Y = 38 else
"110111011111" when X = 58 AND Y = 38 else
"110111011111" when X = 59 AND Y = 38 else
"111111111111" when X = 60 AND Y = 38 else
"111111111111" when X = 61 AND Y = 38 else
"111111111111" when X = 62 AND Y = 38 else
"111111111111" when X = 63 AND Y = 38 else
"111111111111" when X = 64 AND Y = 38 else
"111111111111" when X = 65 AND Y = 38 else
"111111111111" when X = 66 AND Y = 38 else
"111111111111" when X = 67 AND Y = 38 else
"111111111111" when X = 68 AND Y = 38 else
"111111111111" when X = 69 AND Y = 38 else
"111111111111" when X = 70 AND Y = 38 else
"111111111111" when X = 71 AND Y = 38 else
"111111111111" when X = 72 AND Y = 38 else
"111111111111" when X = 73 AND Y = 38 else
"111111111111" when X = 74 AND Y = 38 else
"111111111111" when X = 75 AND Y = 38 else
"111111111111" when X = 76 AND Y = 38 else
"111111111111" when X = 77 AND Y = 38 else
"111111111111" when X = 78 AND Y = 38 else
"111111111111" when X = 79 AND Y = 38 else
"111111111111" when X = 80 AND Y = 38 else
"111111111111" when X = 81 AND Y = 38 else
"111111111111" when X = 82 AND Y = 38 else
"111111111111" when X = 83 AND Y = 38 else
"111111111111" when X = 84 AND Y = 38 else
"111111111111" when X = 85 AND Y = 38 else
"111111111111" when X = 86 AND Y = 38 else
"111111111111" when X = 87 AND Y = 38 else
"111111111111" when X = 88 AND Y = 38 else
"111111111111" when X = 89 AND Y = 38 else
"111111111111" when X = 90 AND Y = 38 else
"111111111111" when X = 91 AND Y = 38 else
"111111111111" when X = 92 AND Y = 38 else
"111111111111" when X = 93 AND Y = 38 else
"111111111111" when X = 94 AND Y = 38 else
"111111111111" when X = 95 AND Y = 38 else
"111111111111" when X = 96 AND Y = 38 else
"111111111111" when X = 97 AND Y = 38 else
"111111111111" when X = 98 AND Y = 38 else
"111111111111" when X = 99 AND Y = 38 else
"111111111111" when X = 100 AND Y = 38 else
"111111111111" when X = 101 AND Y = 38 else
"111111111111" when X = 102 AND Y = 38 else
"111111111111" when X = 103 AND Y = 38 else
"111111111111" when X = 104 AND Y = 38 else
"111111111111" when X = 105 AND Y = 38 else
"111111111111" when X = 106 AND Y = 38 else
"111111111111" when X = 107 AND Y = 38 else
"111111111111" when X = 108 AND Y = 38 else
"111111111111" when X = 109 AND Y = 38 else
"111111111111" when X = 110 AND Y = 38 else
"111111111111" when X = 111 AND Y = 38 else
"111111111111" when X = 112 AND Y = 38 else
"111111111111" when X = 113 AND Y = 38 else
"111111111111" when X = 114 AND Y = 38 else
"111111111111" when X = 115 AND Y = 38 else
"111111111111" when X = 116 AND Y = 38 else
"111111111111" when X = 117 AND Y = 38 else
"111111111111" when X = 118 AND Y = 38 else
"111111111111" when X = 119 AND Y = 38 else
"111111111111" when X = 120 AND Y = 38 else
"111111111111" when X = 121 AND Y = 38 else
"111111111111" when X = 122 AND Y = 38 else
"111111111111" when X = 123 AND Y = 38 else
"111111111111" when X = 124 AND Y = 38 else
"111111111111" when X = 125 AND Y = 38 else
"111111111111" when X = 126 AND Y = 38 else
"111111111111" when X = 127 AND Y = 38 else
"111111111111" when X = 128 AND Y = 38 else
"111111111111" when X = 129 AND Y = 38 else
"111111111111" when X = 130 AND Y = 38 else
"111111111111" when X = 131 AND Y = 38 else
"111111111111" when X = 132 AND Y = 38 else
"111111111111" when X = 133 AND Y = 38 else
"111111111111" when X = 134 AND Y = 38 else
"111111111111" when X = 135 AND Y = 38 else
"111111111111" when X = 136 AND Y = 38 else
"111111111111" when X = 137 AND Y = 38 else
"111111111111" when X = 138 AND Y = 38 else
"111111111111" when X = 139 AND Y = 38 else
"111111111111" when X = 140 AND Y = 38 else
"111111111111" when X = 141 AND Y = 38 else
"111111111111" when X = 142 AND Y = 38 else
"111111111111" when X = 143 AND Y = 38 else
"111111111111" when X = 144 AND Y = 38 else
"111111111111" when X = 145 AND Y = 38 else
"111111111111" when X = 146 AND Y = 38 else
"111111111111" when X = 147 AND Y = 38 else
"111111111111" when X = 148 AND Y = 38 else
"111111111111" when X = 149 AND Y = 38 else
"111111111111" when X = 150 AND Y = 38 else
"111111111111" when X = 151 AND Y = 38 else
"111111111111" when X = 152 AND Y = 38 else
"111111111111" when X = 153 AND Y = 38 else
"111111111111" when X = 154 AND Y = 38 else
"111111111111" when X = 155 AND Y = 38 else
"111111111111" when X = 156 AND Y = 38 else
"111111111111" when X = 157 AND Y = 38 else
"111111111111" when X = 158 AND Y = 38 else
"111111111111" when X = 159 AND Y = 38 else
"111111111111" when X = 160 AND Y = 38 else
"111111111111" when X = 161 AND Y = 38 else
"111111111111" when X = 162 AND Y = 38 else
"111111111111" when X = 163 AND Y = 38 else
"111111111111" when X = 164 AND Y = 38 else
"111111111111" when X = 165 AND Y = 38 else
"111111111111" when X = 166 AND Y = 38 else
"111111111111" when X = 167 AND Y = 38 else
"111111111111" when X = 168 AND Y = 38 else
"111111111111" when X = 169 AND Y = 38 else
"111111111111" when X = 170 AND Y = 38 else
"111111111111" when X = 171 AND Y = 38 else
"111111111111" when X = 172 AND Y = 38 else
"111111111111" when X = 173 AND Y = 38 else
"111111111111" when X = 174 AND Y = 38 else
"111111111111" when X = 175 AND Y = 38 else
"111111111111" when X = 176 AND Y = 38 else
"111111111111" when X = 177 AND Y = 38 else
"111111111111" when X = 178 AND Y = 38 else
"111111111111" when X = 179 AND Y = 38 else
"111111111111" when X = 180 AND Y = 38 else
"111111111111" when X = 181 AND Y = 38 else
"111111111111" when X = 182 AND Y = 38 else
"111111111111" when X = 183 AND Y = 38 else
"111111111111" when X = 184 AND Y = 38 else
"111111111111" when X = 185 AND Y = 38 else
"111111111111" when X = 186 AND Y = 38 else
"111111111111" when X = 187 AND Y = 38 else
"111111111111" when X = 188 AND Y = 38 else
"111111111111" when X = 189 AND Y = 38 else
"111111111111" when X = 190 AND Y = 38 else
"111111111111" when X = 191 AND Y = 38 else
"111111111111" when X = 192 AND Y = 38 else
"111111111111" when X = 193 AND Y = 38 else
"111111111111" when X = 194 AND Y = 38 else
"111111111111" when X = 195 AND Y = 38 else
"111111111111" when X = 196 AND Y = 38 else
"111111111111" when X = 197 AND Y = 38 else
"111111111111" when X = 198 AND Y = 38 else
"111111111111" when X = 199 AND Y = 38 else
"000000000000" when X = 200 AND Y = 38 else
"000000000000" when X = 201 AND Y = 38 else
"000000000000" when X = 202 AND Y = 38 else
"000000000000" when X = 203 AND Y = 38 else
"000000000000" when X = 204 AND Y = 38 else
"000000000000" when X = 205 AND Y = 38 else
"000000000000" when X = 206 AND Y = 38 else
"000000000000" when X = 207 AND Y = 38 else
"000000000000" when X = 208 AND Y = 38 else
"000000000000" when X = 209 AND Y = 38 else
"000000000000" when X = 210 AND Y = 38 else
"000000000000" when X = 211 AND Y = 38 else
"000000000000" when X = 212 AND Y = 38 else
"000000000000" when X = 213 AND Y = 38 else
"000000000000" when X = 214 AND Y = 38 else
"111111111111" when X = 215 AND Y = 38 else
"111111111111" when X = 216 AND Y = 38 else
"111111111111" when X = 217 AND Y = 38 else
"111111111111" when X = 218 AND Y = 38 else
"111111111111" when X = 219 AND Y = 38 else
"111111111111" when X = 220 AND Y = 38 else
"111111111111" when X = 221 AND Y = 38 else
"111111111111" when X = 222 AND Y = 38 else
"111111111111" when X = 223 AND Y = 38 else
"111111111111" when X = 224 AND Y = 38 else
"111111111111" when X = 225 AND Y = 38 else
"111111111111" when X = 226 AND Y = 38 else
"111111111111" when X = 227 AND Y = 38 else
"111111111111" when X = 228 AND Y = 38 else
"111111111111" when X = 229 AND Y = 38 else
"111111111111" when X = 230 AND Y = 38 else
"111111111111" when X = 231 AND Y = 38 else
"111111111111" when X = 232 AND Y = 38 else
"111111111111" when X = 233 AND Y = 38 else
"111111111111" when X = 234 AND Y = 38 else
"111111111111" when X = 235 AND Y = 38 else
"111111111111" when X = 236 AND Y = 38 else
"111111111111" when X = 237 AND Y = 38 else
"111111111111" when X = 238 AND Y = 38 else
"111111111111" when X = 239 AND Y = 38 else
"111111111111" when X = 240 AND Y = 38 else
"111111111111" when X = 241 AND Y = 38 else
"111111111111" when X = 242 AND Y = 38 else
"111111111111" when X = 243 AND Y = 38 else
"111111111111" when X = 244 AND Y = 38 else
"111111111111" when X = 245 AND Y = 38 else
"111111111111" when X = 246 AND Y = 38 else
"111111111111" when X = 247 AND Y = 38 else
"111111111111" when X = 248 AND Y = 38 else
"111111111111" when X = 249 AND Y = 38 else
"111111111111" when X = 250 AND Y = 38 else
"111111111111" when X = 251 AND Y = 38 else
"111111111111" when X = 252 AND Y = 38 else
"111111111111" when X = 253 AND Y = 38 else
"111111111111" when X = 254 AND Y = 38 else
"111111111111" when X = 255 AND Y = 38 else
"111111111111" when X = 256 AND Y = 38 else
"111111111111" when X = 257 AND Y = 38 else
"111111111111" when X = 258 AND Y = 38 else
"111111111111" when X = 259 AND Y = 38 else
"110111011111" when X = 260 AND Y = 38 else
"110111011111" when X = 261 AND Y = 38 else
"110111011111" when X = 262 AND Y = 38 else
"110111011111" when X = 263 AND Y = 38 else
"110111011111" when X = 264 AND Y = 38 else
"110111011111" when X = 265 AND Y = 38 else
"110111011111" when X = 266 AND Y = 38 else
"110111011111" when X = 267 AND Y = 38 else
"110111011111" when X = 268 AND Y = 38 else
"110111011111" when X = 269 AND Y = 38 else
"110111011111" when X = 270 AND Y = 38 else
"110111011111" when X = 271 AND Y = 38 else
"110111011111" when X = 272 AND Y = 38 else
"110111011111" when X = 273 AND Y = 38 else
"110111011111" when X = 274 AND Y = 38 else
"110111011111" when X = 275 AND Y = 38 else
"110111011111" when X = 276 AND Y = 38 else
"110111011111" when X = 277 AND Y = 38 else
"110111011111" when X = 278 AND Y = 38 else
"110111011111" when X = 279 AND Y = 38 else
"000000000000" when X = 280 AND Y = 38 else
"000000000000" when X = 281 AND Y = 38 else
"000000000000" when X = 282 AND Y = 38 else
"000000000000" when X = 283 AND Y = 38 else
"000000000000" when X = 284 AND Y = 38 else
"000000000000" when X = 285 AND Y = 38 else
"000000000000" when X = 286 AND Y = 38 else
"000000000000" when X = 287 AND Y = 38 else
"000000000000" when X = 288 AND Y = 38 else
"000000000000" when X = 289 AND Y = 38 else
"000000000000" when X = 290 AND Y = 38 else
"000000000000" when X = 291 AND Y = 38 else
"000000000000" when X = 292 AND Y = 38 else
"000000000000" when X = 293 AND Y = 38 else
"000000000000" when X = 294 AND Y = 38 else
"000000000000" when X = 295 AND Y = 38 else
"000000000000" when X = 296 AND Y = 38 else
"000000000000" when X = 297 AND Y = 38 else
"000000000000" when X = 298 AND Y = 38 else
"000000000000" when X = 299 AND Y = 38 else
"000000000000" when X = 300 AND Y = 38 else
"000000000000" when X = 301 AND Y = 38 else
"000000000000" when X = 302 AND Y = 38 else
"000000000000" when X = 303 AND Y = 38 else
"000000000000" when X = 304 AND Y = 38 else
"000000000000" when X = 305 AND Y = 38 else
"000000000000" when X = 306 AND Y = 38 else
"000000000000" when X = 307 AND Y = 38 else
"000000000000" when X = 308 AND Y = 38 else
"000000000000" when X = 309 AND Y = 38 else
"000000000000" when X = 310 AND Y = 38 else
"000000000000" when X = 311 AND Y = 38 else
"000000000000" when X = 312 AND Y = 38 else
"000000000000" when X = 313 AND Y = 38 else
"000000000000" when X = 314 AND Y = 38 else
"000000000000" when X = 315 AND Y = 38 else
"000000000000" when X = 316 AND Y = 38 else
"000000000000" when X = 317 AND Y = 38 else
"000000000000" when X = 318 AND Y = 38 else
"000000000000" when X = 319 AND Y = 38 else
"000000000000" when X = 320 AND Y = 38 else
"000000000000" when X = 321 AND Y = 38 else
"000000000000" when X = 322 AND Y = 38 else
"000000000000" when X = 323 AND Y = 38 else
"000000000000" when X = 324 AND Y = 38 else
"000000000000" when X = 0 AND Y = 39 else
"000000000000" when X = 1 AND Y = 39 else
"000000000000" when X = 2 AND Y = 39 else
"000000000000" when X = 3 AND Y = 39 else
"000000000000" when X = 4 AND Y = 39 else
"000000000000" when X = 5 AND Y = 39 else
"000000000000" when X = 6 AND Y = 39 else
"000000000000" when X = 7 AND Y = 39 else
"000000000000" when X = 8 AND Y = 39 else
"000000000000" when X = 9 AND Y = 39 else
"000000000000" when X = 10 AND Y = 39 else
"000000000000" when X = 11 AND Y = 39 else
"000000000000" when X = 12 AND Y = 39 else
"000000000000" when X = 13 AND Y = 39 else
"000000000000" when X = 14 AND Y = 39 else
"000000000000" when X = 15 AND Y = 39 else
"000000000000" when X = 16 AND Y = 39 else
"000000000000" when X = 17 AND Y = 39 else
"000000000000" when X = 18 AND Y = 39 else
"000000000000" when X = 19 AND Y = 39 else
"000000000000" when X = 20 AND Y = 39 else
"000000000000" when X = 21 AND Y = 39 else
"000000000000" when X = 22 AND Y = 39 else
"000000000000" when X = 23 AND Y = 39 else
"000000000000" when X = 24 AND Y = 39 else
"000000000000" when X = 25 AND Y = 39 else
"000000000000" when X = 26 AND Y = 39 else
"000000000000" when X = 27 AND Y = 39 else
"000000000000" when X = 28 AND Y = 39 else
"000000000000" when X = 29 AND Y = 39 else
"000000000000" when X = 30 AND Y = 39 else
"000000000000" when X = 31 AND Y = 39 else
"000000000000" when X = 32 AND Y = 39 else
"000000000000" when X = 33 AND Y = 39 else
"000000000000" when X = 34 AND Y = 39 else
"000000000000" when X = 35 AND Y = 39 else
"000000000000" when X = 36 AND Y = 39 else
"000000000000" when X = 37 AND Y = 39 else
"000000000000" when X = 38 AND Y = 39 else
"000000000000" when X = 39 AND Y = 39 else
"100010011101" when X = 40 AND Y = 39 else
"100010011101" when X = 41 AND Y = 39 else
"100010011101" when X = 42 AND Y = 39 else
"100010011101" when X = 43 AND Y = 39 else
"100010011101" when X = 44 AND Y = 39 else
"100010011101" when X = 45 AND Y = 39 else
"100010011101" when X = 46 AND Y = 39 else
"100010011101" when X = 47 AND Y = 39 else
"100010011101" when X = 48 AND Y = 39 else
"100010011101" when X = 49 AND Y = 39 else
"110111011111" when X = 50 AND Y = 39 else
"110111011111" when X = 51 AND Y = 39 else
"110111011111" when X = 52 AND Y = 39 else
"110111011111" when X = 53 AND Y = 39 else
"110111011111" when X = 54 AND Y = 39 else
"110111011111" when X = 55 AND Y = 39 else
"110111011111" when X = 56 AND Y = 39 else
"110111011111" when X = 57 AND Y = 39 else
"110111011111" when X = 58 AND Y = 39 else
"110111011111" when X = 59 AND Y = 39 else
"111111111111" when X = 60 AND Y = 39 else
"111111111111" when X = 61 AND Y = 39 else
"111111111111" when X = 62 AND Y = 39 else
"111111111111" when X = 63 AND Y = 39 else
"111111111111" when X = 64 AND Y = 39 else
"111111111111" when X = 65 AND Y = 39 else
"111111111111" when X = 66 AND Y = 39 else
"111111111111" when X = 67 AND Y = 39 else
"111111111111" when X = 68 AND Y = 39 else
"111111111111" when X = 69 AND Y = 39 else
"111111111111" when X = 70 AND Y = 39 else
"111111111111" when X = 71 AND Y = 39 else
"111111111111" when X = 72 AND Y = 39 else
"111111111111" when X = 73 AND Y = 39 else
"111111111111" when X = 74 AND Y = 39 else
"111111111111" when X = 75 AND Y = 39 else
"111111111111" when X = 76 AND Y = 39 else
"111111111111" when X = 77 AND Y = 39 else
"111111111111" when X = 78 AND Y = 39 else
"111111111111" when X = 79 AND Y = 39 else
"111111111111" when X = 80 AND Y = 39 else
"111111111111" when X = 81 AND Y = 39 else
"111111111111" when X = 82 AND Y = 39 else
"111111111111" when X = 83 AND Y = 39 else
"111111111111" when X = 84 AND Y = 39 else
"111111111111" when X = 85 AND Y = 39 else
"111111111111" when X = 86 AND Y = 39 else
"111111111111" when X = 87 AND Y = 39 else
"111111111111" when X = 88 AND Y = 39 else
"111111111111" when X = 89 AND Y = 39 else
"111111111111" when X = 90 AND Y = 39 else
"111111111111" when X = 91 AND Y = 39 else
"111111111111" when X = 92 AND Y = 39 else
"111111111111" when X = 93 AND Y = 39 else
"111111111111" when X = 94 AND Y = 39 else
"111111111111" when X = 95 AND Y = 39 else
"111111111111" when X = 96 AND Y = 39 else
"111111111111" when X = 97 AND Y = 39 else
"111111111111" when X = 98 AND Y = 39 else
"111111111111" when X = 99 AND Y = 39 else
"111111111111" when X = 100 AND Y = 39 else
"111111111111" when X = 101 AND Y = 39 else
"111111111111" when X = 102 AND Y = 39 else
"111111111111" when X = 103 AND Y = 39 else
"111111111111" when X = 104 AND Y = 39 else
"111111111111" when X = 105 AND Y = 39 else
"111111111111" when X = 106 AND Y = 39 else
"111111111111" when X = 107 AND Y = 39 else
"111111111111" when X = 108 AND Y = 39 else
"111111111111" when X = 109 AND Y = 39 else
"111111111111" when X = 110 AND Y = 39 else
"111111111111" when X = 111 AND Y = 39 else
"111111111111" when X = 112 AND Y = 39 else
"111111111111" when X = 113 AND Y = 39 else
"111111111111" when X = 114 AND Y = 39 else
"111111111111" when X = 115 AND Y = 39 else
"111111111111" when X = 116 AND Y = 39 else
"111111111111" when X = 117 AND Y = 39 else
"111111111111" when X = 118 AND Y = 39 else
"111111111111" when X = 119 AND Y = 39 else
"111111111111" when X = 120 AND Y = 39 else
"111111111111" when X = 121 AND Y = 39 else
"111111111111" when X = 122 AND Y = 39 else
"111111111111" when X = 123 AND Y = 39 else
"111111111111" when X = 124 AND Y = 39 else
"111111111111" when X = 125 AND Y = 39 else
"111111111111" when X = 126 AND Y = 39 else
"111111111111" when X = 127 AND Y = 39 else
"111111111111" when X = 128 AND Y = 39 else
"111111111111" when X = 129 AND Y = 39 else
"111111111111" when X = 130 AND Y = 39 else
"111111111111" when X = 131 AND Y = 39 else
"111111111111" when X = 132 AND Y = 39 else
"111111111111" when X = 133 AND Y = 39 else
"111111111111" when X = 134 AND Y = 39 else
"111111111111" when X = 135 AND Y = 39 else
"111111111111" when X = 136 AND Y = 39 else
"111111111111" when X = 137 AND Y = 39 else
"111111111111" when X = 138 AND Y = 39 else
"111111111111" when X = 139 AND Y = 39 else
"111111111111" when X = 140 AND Y = 39 else
"111111111111" when X = 141 AND Y = 39 else
"111111111111" when X = 142 AND Y = 39 else
"111111111111" when X = 143 AND Y = 39 else
"111111111111" when X = 144 AND Y = 39 else
"111111111111" when X = 145 AND Y = 39 else
"111111111111" when X = 146 AND Y = 39 else
"111111111111" when X = 147 AND Y = 39 else
"111111111111" when X = 148 AND Y = 39 else
"111111111111" when X = 149 AND Y = 39 else
"111111111111" when X = 150 AND Y = 39 else
"111111111111" when X = 151 AND Y = 39 else
"111111111111" when X = 152 AND Y = 39 else
"111111111111" when X = 153 AND Y = 39 else
"111111111111" when X = 154 AND Y = 39 else
"111111111111" when X = 155 AND Y = 39 else
"111111111111" when X = 156 AND Y = 39 else
"111111111111" when X = 157 AND Y = 39 else
"111111111111" when X = 158 AND Y = 39 else
"111111111111" when X = 159 AND Y = 39 else
"111111111111" when X = 160 AND Y = 39 else
"111111111111" when X = 161 AND Y = 39 else
"111111111111" when X = 162 AND Y = 39 else
"111111111111" when X = 163 AND Y = 39 else
"111111111111" when X = 164 AND Y = 39 else
"111111111111" when X = 165 AND Y = 39 else
"111111111111" when X = 166 AND Y = 39 else
"111111111111" when X = 167 AND Y = 39 else
"111111111111" when X = 168 AND Y = 39 else
"111111111111" when X = 169 AND Y = 39 else
"111111111111" when X = 170 AND Y = 39 else
"111111111111" when X = 171 AND Y = 39 else
"111111111111" when X = 172 AND Y = 39 else
"111111111111" when X = 173 AND Y = 39 else
"111111111111" when X = 174 AND Y = 39 else
"111111111111" when X = 175 AND Y = 39 else
"111111111111" when X = 176 AND Y = 39 else
"111111111111" when X = 177 AND Y = 39 else
"111111111111" when X = 178 AND Y = 39 else
"111111111111" when X = 179 AND Y = 39 else
"111111111111" when X = 180 AND Y = 39 else
"111111111111" when X = 181 AND Y = 39 else
"111111111111" when X = 182 AND Y = 39 else
"111111111111" when X = 183 AND Y = 39 else
"111111111111" when X = 184 AND Y = 39 else
"111111111111" when X = 185 AND Y = 39 else
"111111111111" when X = 186 AND Y = 39 else
"111111111111" when X = 187 AND Y = 39 else
"111111111111" when X = 188 AND Y = 39 else
"111111111111" when X = 189 AND Y = 39 else
"111111111111" when X = 190 AND Y = 39 else
"111111111111" when X = 191 AND Y = 39 else
"111111111111" when X = 192 AND Y = 39 else
"111111111111" when X = 193 AND Y = 39 else
"111111111111" when X = 194 AND Y = 39 else
"111111111111" when X = 195 AND Y = 39 else
"111111111111" when X = 196 AND Y = 39 else
"111111111111" when X = 197 AND Y = 39 else
"111111111111" when X = 198 AND Y = 39 else
"111111111111" when X = 199 AND Y = 39 else
"000000000000" when X = 200 AND Y = 39 else
"000000000000" when X = 201 AND Y = 39 else
"000000000000" when X = 202 AND Y = 39 else
"000000000000" when X = 203 AND Y = 39 else
"000000000000" when X = 204 AND Y = 39 else
"000000000000" when X = 205 AND Y = 39 else
"000000000000" when X = 206 AND Y = 39 else
"000000000000" when X = 207 AND Y = 39 else
"000000000000" when X = 208 AND Y = 39 else
"000000000000" when X = 209 AND Y = 39 else
"000000000000" when X = 210 AND Y = 39 else
"000000000000" when X = 211 AND Y = 39 else
"000000000000" when X = 212 AND Y = 39 else
"000000000000" when X = 213 AND Y = 39 else
"000000000000" when X = 214 AND Y = 39 else
"111111111111" when X = 215 AND Y = 39 else
"111111111111" when X = 216 AND Y = 39 else
"111111111111" when X = 217 AND Y = 39 else
"111111111111" when X = 218 AND Y = 39 else
"111111111111" when X = 219 AND Y = 39 else
"111111111111" when X = 220 AND Y = 39 else
"111111111111" when X = 221 AND Y = 39 else
"111111111111" when X = 222 AND Y = 39 else
"111111111111" when X = 223 AND Y = 39 else
"111111111111" when X = 224 AND Y = 39 else
"111111111111" when X = 225 AND Y = 39 else
"111111111111" when X = 226 AND Y = 39 else
"111111111111" when X = 227 AND Y = 39 else
"111111111111" when X = 228 AND Y = 39 else
"111111111111" when X = 229 AND Y = 39 else
"111111111111" when X = 230 AND Y = 39 else
"111111111111" when X = 231 AND Y = 39 else
"111111111111" when X = 232 AND Y = 39 else
"111111111111" when X = 233 AND Y = 39 else
"111111111111" when X = 234 AND Y = 39 else
"111111111111" when X = 235 AND Y = 39 else
"111111111111" when X = 236 AND Y = 39 else
"111111111111" when X = 237 AND Y = 39 else
"111111111111" when X = 238 AND Y = 39 else
"111111111111" when X = 239 AND Y = 39 else
"111111111111" when X = 240 AND Y = 39 else
"111111111111" when X = 241 AND Y = 39 else
"111111111111" when X = 242 AND Y = 39 else
"111111111111" when X = 243 AND Y = 39 else
"111111111111" when X = 244 AND Y = 39 else
"111111111111" when X = 245 AND Y = 39 else
"111111111111" when X = 246 AND Y = 39 else
"111111111111" when X = 247 AND Y = 39 else
"111111111111" when X = 248 AND Y = 39 else
"111111111111" when X = 249 AND Y = 39 else
"111111111111" when X = 250 AND Y = 39 else
"111111111111" when X = 251 AND Y = 39 else
"111111111111" when X = 252 AND Y = 39 else
"111111111111" when X = 253 AND Y = 39 else
"111111111111" when X = 254 AND Y = 39 else
"111111111111" when X = 255 AND Y = 39 else
"111111111111" when X = 256 AND Y = 39 else
"111111111111" when X = 257 AND Y = 39 else
"111111111111" when X = 258 AND Y = 39 else
"111111111111" when X = 259 AND Y = 39 else
"110111011111" when X = 260 AND Y = 39 else
"110111011111" when X = 261 AND Y = 39 else
"110111011111" when X = 262 AND Y = 39 else
"110111011111" when X = 263 AND Y = 39 else
"110111011111" when X = 264 AND Y = 39 else
"110111011111" when X = 265 AND Y = 39 else
"110111011111" when X = 266 AND Y = 39 else
"110111011111" when X = 267 AND Y = 39 else
"110111011111" when X = 268 AND Y = 39 else
"110111011111" when X = 269 AND Y = 39 else
"110111011111" when X = 270 AND Y = 39 else
"110111011111" when X = 271 AND Y = 39 else
"110111011111" when X = 272 AND Y = 39 else
"110111011111" when X = 273 AND Y = 39 else
"110111011111" when X = 274 AND Y = 39 else
"110111011111" when X = 275 AND Y = 39 else
"110111011111" when X = 276 AND Y = 39 else
"110111011111" when X = 277 AND Y = 39 else
"110111011111" when X = 278 AND Y = 39 else
"110111011111" when X = 279 AND Y = 39 else
"000000000000" when X = 280 AND Y = 39 else
"000000000000" when X = 281 AND Y = 39 else
"000000000000" when X = 282 AND Y = 39 else
"000000000000" when X = 283 AND Y = 39 else
"000000000000" when X = 284 AND Y = 39 else
"000000000000" when X = 285 AND Y = 39 else
"000000000000" when X = 286 AND Y = 39 else
"000000000000" when X = 287 AND Y = 39 else
"000000000000" when X = 288 AND Y = 39 else
"000000000000" when X = 289 AND Y = 39 else
"000000000000" when X = 290 AND Y = 39 else
"000000000000" when X = 291 AND Y = 39 else
"000000000000" when X = 292 AND Y = 39 else
"000000000000" when X = 293 AND Y = 39 else
"000000000000" when X = 294 AND Y = 39 else
"000000000000" when X = 295 AND Y = 39 else
"000000000000" when X = 296 AND Y = 39 else
"000000000000" when X = 297 AND Y = 39 else
"000000000000" when X = 298 AND Y = 39 else
"000000000000" when X = 299 AND Y = 39 else
"000000000000" when X = 300 AND Y = 39 else
"000000000000" when X = 301 AND Y = 39 else
"000000000000" when X = 302 AND Y = 39 else
"000000000000" when X = 303 AND Y = 39 else
"000000000000" when X = 304 AND Y = 39 else
"000000000000" when X = 305 AND Y = 39 else
"000000000000" when X = 306 AND Y = 39 else
"000000000000" when X = 307 AND Y = 39 else
"000000000000" when X = 308 AND Y = 39 else
"000000000000" when X = 309 AND Y = 39 else
"000000000000" when X = 310 AND Y = 39 else
"000000000000" when X = 311 AND Y = 39 else
"000000000000" when X = 312 AND Y = 39 else
"000000000000" when X = 313 AND Y = 39 else
"000000000000" when X = 314 AND Y = 39 else
"000000000000" when X = 315 AND Y = 39 else
"000000000000" when X = 316 AND Y = 39 else
"000000000000" when X = 317 AND Y = 39 else
"000000000000" when X = 318 AND Y = 39 else
"000000000000" when X = 319 AND Y = 39 else
"000000000000" when X = 320 AND Y = 39 else
"000000000000" when X = 321 AND Y = 39 else
"000000000000" when X = 322 AND Y = 39 else
"000000000000" when X = 323 AND Y = 39 else
"000000000000" when X = 324 AND Y = 39 else
"000000000000" when X = 0 AND Y = 40 else
"000000000000" when X = 1 AND Y = 40 else
"000000000000" when X = 2 AND Y = 40 else
"000000000000" when X = 3 AND Y = 40 else
"000000000000" when X = 4 AND Y = 40 else
"000000000000" when X = 5 AND Y = 40 else
"000000000000" when X = 6 AND Y = 40 else
"000000000000" when X = 7 AND Y = 40 else
"000000000000" when X = 8 AND Y = 40 else
"000000000000" when X = 9 AND Y = 40 else
"000000000000" when X = 10 AND Y = 40 else
"000000000000" when X = 11 AND Y = 40 else
"000000000000" when X = 12 AND Y = 40 else
"000000000000" when X = 13 AND Y = 40 else
"000000000000" when X = 14 AND Y = 40 else
"000000000000" when X = 15 AND Y = 40 else
"000000000000" when X = 16 AND Y = 40 else
"000000000000" when X = 17 AND Y = 40 else
"000000000000" when X = 18 AND Y = 40 else
"000000000000" when X = 19 AND Y = 40 else
"000000000000" when X = 20 AND Y = 40 else
"000000000000" when X = 21 AND Y = 40 else
"000000000000" when X = 22 AND Y = 40 else
"000000000000" when X = 23 AND Y = 40 else
"000000000000" when X = 24 AND Y = 40 else
"000000000000" when X = 25 AND Y = 40 else
"000000000000" when X = 26 AND Y = 40 else
"000000000000" when X = 27 AND Y = 40 else
"000000000000" when X = 28 AND Y = 40 else
"000000000000" when X = 29 AND Y = 40 else
"000000000000" when X = 30 AND Y = 40 else
"000000000000" when X = 31 AND Y = 40 else
"000000000000" when X = 32 AND Y = 40 else
"000000000000" when X = 33 AND Y = 40 else
"000000000000" when X = 34 AND Y = 40 else
"000000000000" when X = 35 AND Y = 40 else
"000000000000" when X = 36 AND Y = 40 else
"000000000000" when X = 37 AND Y = 40 else
"000000000000" when X = 38 AND Y = 40 else
"000000000000" when X = 39 AND Y = 40 else
"100010011101" when X = 40 AND Y = 40 else
"100010011101" when X = 41 AND Y = 40 else
"100010011101" when X = 42 AND Y = 40 else
"100010011101" when X = 43 AND Y = 40 else
"100010011101" when X = 44 AND Y = 40 else
"100010011101" when X = 45 AND Y = 40 else
"100010011101" when X = 46 AND Y = 40 else
"100010011101" when X = 47 AND Y = 40 else
"100010011101" when X = 48 AND Y = 40 else
"100010011101" when X = 49 AND Y = 40 else
"110111011111" when X = 50 AND Y = 40 else
"110111011111" when X = 51 AND Y = 40 else
"110111011111" when X = 52 AND Y = 40 else
"110111011111" when X = 53 AND Y = 40 else
"110111011111" when X = 54 AND Y = 40 else
"110111011111" when X = 55 AND Y = 40 else
"110111011111" when X = 56 AND Y = 40 else
"110111011111" when X = 57 AND Y = 40 else
"110111011111" when X = 58 AND Y = 40 else
"110111011111" when X = 59 AND Y = 40 else
"111111111111" when X = 60 AND Y = 40 else
"111111111111" when X = 61 AND Y = 40 else
"111111111111" when X = 62 AND Y = 40 else
"111111111111" when X = 63 AND Y = 40 else
"111111111111" when X = 64 AND Y = 40 else
"111111111111" when X = 65 AND Y = 40 else
"111111111111" when X = 66 AND Y = 40 else
"111111111111" when X = 67 AND Y = 40 else
"111111111111" when X = 68 AND Y = 40 else
"111111111111" when X = 69 AND Y = 40 else
"111111111111" when X = 70 AND Y = 40 else
"111111111111" when X = 71 AND Y = 40 else
"111111111111" when X = 72 AND Y = 40 else
"111111111111" when X = 73 AND Y = 40 else
"111111111111" when X = 74 AND Y = 40 else
"111111111111" when X = 75 AND Y = 40 else
"111111111111" when X = 76 AND Y = 40 else
"111111111111" when X = 77 AND Y = 40 else
"111111111111" when X = 78 AND Y = 40 else
"111111111111" when X = 79 AND Y = 40 else
"111111111111" when X = 80 AND Y = 40 else
"111111111111" when X = 81 AND Y = 40 else
"111111111111" when X = 82 AND Y = 40 else
"111111111111" when X = 83 AND Y = 40 else
"111111111111" when X = 84 AND Y = 40 else
"111111111111" when X = 85 AND Y = 40 else
"111111111111" when X = 86 AND Y = 40 else
"111111111111" when X = 87 AND Y = 40 else
"111111111111" when X = 88 AND Y = 40 else
"111111111111" when X = 89 AND Y = 40 else
"111111111111" when X = 90 AND Y = 40 else
"111111111111" when X = 91 AND Y = 40 else
"111111111111" when X = 92 AND Y = 40 else
"111111111111" when X = 93 AND Y = 40 else
"111111111111" when X = 94 AND Y = 40 else
"111111111111" when X = 95 AND Y = 40 else
"111111111111" when X = 96 AND Y = 40 else
"111111111111" when X = 97 AND Y = 40 else
"111111111111" when X = 98 AND Y = 40 else
"111111111111" when X = 99 AND Y = 40 else
"111111111111" when X = 100 AND Y = 40 else
"111111111111" when X = 101 AND Y = 40 else
"111111111111" when X = 102 AND Y = 40 else
"111111111111" when X = 103 AND Y = 40 else
"111111111111" when X = 104 AND Y = 40 else
"111111111111" when X = 105 AND Y = 40 else
"111111111111" when X = 106 AND Y = 40 else
"111111111111" when X = 107 AND Y = 40 else
"111111111111" when X = 108 AND Y = 40 else
"111111111111" when X = 109 AND Y = 40 else
"111111111111" when X = 110 AND Y = 40 else
"111111111111" when X = 111 AND Y = 40 else
"111111111111" when X = 112 AND Y = 40 else
"111111111111" when X = 113 AND Y = 40 else
"111111111111" when X = 114 AND Y = 40 else
"111111111111" when X = 115 AND Y = 40 else
"111111111111" when X = 116 AND Y = 40 else
"111111111111" when X = 117 AND Y = 40 else
"111111111111" when X = 118 AND Y = 40 else
"111111111111" when X = 119 AND Y = 40 else
"111111111111" when X = 120 AND Y = 40 else
"111111111111" when X = 121 AND Y = 40 else
"111111111111" when X = 122 AND Y = 40 else
"111111111111" when X = 123 AND Y = 40 else
"111111111111" when X = 124 AND Y = 40 else
"111111111111" when X = 125 AND Y = 40 else
"111111111111" when X = 126 AND Y = 40 else
"111111111111" when X = 127 AND Y = 40 else
"111111111111" when X = 128 AND Y = 40 else
"111111111111" when X = 129 AND Y = 40 else
"111111111111" when X = 130 AND Y = 40 else
"111111111111" when X = 131 AND Y = 40 else
"111111111111" when X = 132 AND Y = 40 else
"111111111111" when X = 133 AND Y = 40 else
"111111111111" when X = 134 AND Y = 40 else
"111111111111" when X = 135 AND Y = 40 else
"111111111111" when X = 136 AND Y = 40 else
"111111111111" when X = 137 AND Y = 40 else
"111111111111" when X = 138 AND Y = 40 else
"111111111111" when X = 139 AND Y = 40 else
"111111111111" when X = 140 AND Y = 40 else
"111111111111" when X = 141 AND Y = 40 else
"111111111111" when X = 142 AND Y = 40 else
"111111111111" when X = 143 AND Y = 40 else
"111111111111" when X = 144 AND Y = 40 else
"111111111111" when X = 145 AND Y = 40 else
"111111111111" when X = 146 AND Y = 40 else
"111111111111" when X = 147 AND Y = 40 else
"111111111111" when X = 148 AND Y = 40 else
"111111111111" when X = 149 AND Y = 40 else
"111111111111" when X = 150 AND Y = 40 else
"111111111111" when X = 151 AND Y = 40 else
"111111111111" when X = 152 AND Y = 40 else
"111111111111" when X = 153 AND Y = 40 else
"111111111111" when X = 154 AND Y = 40 else
"111111111111" when X = 155 AND Y = 40 else
"111111111111" when X = 156 AND Y = 40 else
"111111111111" when X = 157 AND Y = 40 else
"111111111111" when X = 158 AND Y = 40 else
"111111111111" when X = 159 AND Y = 40 else
"111111111111" when X = 160 AND Y = 40 else
"111111111111" when X = 161 AND Y = 40 else
"111111111111" when X = 162 AND Y = 40 else
"111111111111" when X = 163 AND Y = 40 else
"111111111111" when X = 164 AND Y = 40 else
"111111111111" when X = 165 AND Y = 40 else
"111111111111" when X = 166 AND Y = 40 else
"111111111111" when X = 167 AND Y = 40 else
"111111111111" when X = 168 AND Y = 40 else
"111111111111" when X = 169 AND Y = 40 else
"111111111111" when X = 170 AND Y = 40 else
"111111111111" when X = 171 AND Y = 40 else
"111111111111" when X = 172 AND Y = 40 else
"111111111111" when X = 173 AND Y = 40 else
"111111111111" when X = 174 AND Y = 40 else
"111111111111" when X = 175 AND Y = 40 else
"111111111111" when X = 176 AND Y = 40 else
"111111111111" when X = 177 AND Y = 40 else
"111111111111" when X = 178 AND Y = 40 else
"111111111111" when X = 179 AND Y = 40 else
"111111111111" when X = 180 AND Y = 40 else
"111111111111" when X = 181 AND Y = 40 else
"111111111111" when X = 182 AND Y = 40 else
"111111111111" when X = 183 AND Y = 40 else
"111111111111" when X = 184 AND Y = 40 else
"111111111111" when X = 185 AND Y = 40 else
"111111111111" when X = 186 AND Y = 40 else
"111111111111" when X = 187 AND Y = 40 else
"111111111111" when X = 188 AND Y = 40 else
"111111111111" when X = 189 AND Y = 40 else
"111111111111" when X = 190 AND Y = 40 else
"111111111111" when X = 191 AND Y = 40 else
"111111111111" when X = 192 AND Y = 40 else
"111111111111" when X = 193 AND Y = 40 else
"111111111111" when X = 194 AND Y = 40 else
"111111111111" when X = 195 AND Y = 40 else
"111111111111" when X = 196 AND Y = 40 else
"111111111111" when X = 197 AND Y = 40 else
"111111111111" when X = 198 AND Y = 40 else
"111111111111" when X = 199 AND Y = 40 else
"111111111111" when X = 200 AND Y = 40 else
"111111111111" when X = 201 AND Y = 40 else
"111111111111" when X = 202 AND Y = 40 else
"111111111111" when X = 203 AND Y = 40 else
"111111111111" when X = 204 AND Y = 40 else
"111111111111" when X = 205 AND Y = 40 else
"111111111111" when X = 206 AND Y = 40 else
"111111111111" when X = 207 AND Y = 40 else
"111111111111" when X = 208 AND Y = 40 else
"111111111111" when X = 209 AND Y = 40 else
"111111111111" when X = 210 AND Y = 40 else
"111111111111" when X = 211 AND Y = 40 else
"111111111111" when X = 212 AND Y = 40 else
"111111111111" when X = 213 AND Y = 40 else
"111111111111" when X = 214 AND Y = 40 else
"111111111111" when X = 215 AND Y = 40 else
"111111111111" when X = 216 AND Y = 40 else
"111111111111" when X = 217 AND Y = 40 else
"111111111111" when X = 218 AND Y = 40 else
"111111111111" when X = 219 AND Y = 40 else
"111111111111" when X = 220 AND Y = 40 else
"111111111111" when X = 221 AND Y = 40 else
"111111111111" when X = 222 AND Y = 40 else
"111111111111" when X = 223 AND Y = 40 else
"111111111111" when X = 224 AND Y = 40 else
"111111111111" when X = 225 AND Y = 40 else
"111111111111" when X = 226 AND Y = 40 else
"111111111111" when X = 227 AND Y = 40 else
"111111111111" when X = 228 AND Y = 40 else
"111111111111" when X = 229 AND Y = 40 else
"111111111111" when X = 230 AND Y = 40 else
"111111111111" when X = 231 AND Y = 40 else
"111111111111" when X = 232 AND Y = 40 else
"111111111111" when X = 233 AND Y = 40 else
"111111111111" when X = 234 AND Y = 40 else
"111111111111" when X = 235 AND Y = 40 else
"111111111111" when X = 236 AND Y = 40 else
"111111111111" when X = 237 AND Y = 40 else
"111111111111" when X = 238 AND Y = 40 else
"111111111111" when X = 239 AND Y = 40 else
"111111111111" when X = 240 AND Y = 40 else
"111111111111" when X = 241 AND Y = 40 else
"111111111111" when X = 242 AND Y = 40 else
"111111111111" when X = 243 AND Y = 40 else
"111111111111" when X = 244 AND Y = 40 else
"111111111111" when X = 245 AND Y = 40 else
"111111111111" when X = 246 AND Y = 40 else
"111111111111" when X = 247 AND Y = 40 else
"111111111111" when X = 248 AND Y = 40 else
"111111111111" when X = 249 AND Y = 40 else
"111111111111" when X = 250 AND Y = 40 else
"111111111111" when X = 251 AND Y = 40 else
"111111111111" when X = 252 AND Y = 40 else
"111111111111" when X = 253 AND Y = 40 else
"111111111111" when X = 254 AND Y = 40 else
"111111111111" when X = 255 AND Y = 40 else
"111111111111" when X = 256 AND Y = 40 else
"111111111111" when X = 257 AND Y = 40 else
"111111111111" when X = 258 AND Y = 40 else
"111111111111" when X = 259 AND Y = 40 else
"111111111111" when X = 260 AND Y = 40 else
"111111111111" when X = 261 AND Y = 40 else
"111111111111" when X = 262 AND Y = 40 else
"111111111111" when X = 263 AND Y = 40 else
"111111111111" when X = 264 AND Y = 40 else
"110111011111" when X = 265 AND Y = 40 else
"110111011111" when X = 266 AND Y = 40 else
"110111011111" when X = 267 AND Y = 40 else
"110111011111" when X = 268 AND Y = 40 else
"110111011111" when X = 269 AND Y = 40 else
"110111011111" when X = 270 AND Y = 40 else
"110111011111" when X = 271 AND Y = 40 else
"110111011111" when X = 272 AND Y = 40 else
"110111011111" when X = 273 AND Y = 40 else
"110111011111" when X = 274 AND Y = 40 else
"110111011111" when X = 275 AND Y = 40 else
"110111011111" when X = 276 AND Y = 40 else
"110111011111" when X = 277 AND Y = 40 else
"110111011111" when X = 278 AND Y = 40 else
"110111011111" when X = 279 AND Y = 40 else
"000000000000" when X = 280 AND Y = 40 else
"000000000000" when X = 281 AND Y = 40 else
"000000000000" when X = 282 AND Y = 40 else
"000000000000" when X = 283 AND Y = 40 else
"000000000000" when X = 284 AND Y = 40 else
"000000000000" when X = 285 AND Y = 40 else
"000000000000" when X = 286 AND Y = 40 else
"000000000000" when X = 287 AND Y = 40 else
"000000000000" when X = 288 AND Y = 40 else
"000000000000" when X = 289 AND Y = 40 else
"000000000000" when X = 290 AND Y = 40 else
"000000000000" when X = 291 AND Y = 40 else
"000000000000" when X = 292 AND Y = 40 else
"000000000000" when X = 293 AND Y = 40 else
"000000000000" when X = 294 AND Y = 40 else
"000000000000" when X = 295 AND Y = 40 else
"000000000000" when X = 296 AND Y = 40 else
"000000000000" when X = 297 AND Y = 40 else
"000000000000" when X = 298 AND Y = 40 else
"000000000000" when X = 299 AND Y = 40 else
"000000000000" when X = 300 AND Y = 40 else
"000000000000" when X = 301 AND Y = 40 else
"000000000000" when X = 302 AND Y = 40 else
"000000000000" when X = 303 AND Y = 40 else
"000000000000" when X = 304 AND Y = 40 else
"000000000000" when X = 305 AND Y = 40 else
"000000000000" when X = 306 AND Y = 40 else
"000000000000" when X = 307 AND Y = 40 else
"000000000000" when X = 308 AND Y = 40 else
"000000000000" when X = 309 AND Y = 40 else
"000000000000" when X = 310 AND Y = 40 else
"000000000000" when X = 311 AND Y = 40 else
"000000000000" when X = 312 AND Y = 40 else
"000000000000" when X = 313 AND Y = 40 else
"000000000000" when X = 314 AND Y = 40 else
"000000000000" when X = 315 AND Y = 40 else
"000000000000" when X = 316 AND Y = 40 else
"000000000000" when X = 317 AND Y = 40 else
"000000000000" when X = 318 AND Y = 40 else
"000000000000" when X = 319 AND Y = 40 else
"000000000000" when X = 320 AND Y = 40 else
"000000000000" when X = 321 AND Y = 40 else
"000000000000" when X = 322 AND Y = 40 else
"000000000000" when X = 323 AND Y = 40 else
"000000000000" when X = 324 AND Y = 40 else
"000000000000" when X = 0 AND Y = 41 else
"000000000000" when X = 1 AND Y = 41 else
"000000000000" when X = 2 AND Y = 41 else
"000000000000" when X = 3 AND Y = 41 else
"000000000000" when X = 4 AND Y = 41 else
"000000000000" when X = 5 AND Y = 41 else
"000000000000" when X = 6 AND Y = 41 else
"000000000000" when X = 7 AND Y = 41 else
"000000000000" when X = 8 AND Y = 41 else
"000000000000" when X = 9 AND Y = 41 else
"000000000000" when X = 10 AND Y = 41 else
"000000000000" when X = 11 AND Y = 41 else
"000000000000" when X = 12 AND Y = 41 else
"000000000000" when X = 13 AND Y = 41 else
"000000000000" when X = 14 AND Y = 41 else
"000000000000" when X = 15 AND Y = 41 else
"000000000000" when X = 16 AND Y = 41 else
"000000000000" when X = 17 AND Y = 41 else
"000000000000" when X = 18 AND Y = 41 else
"000000000000" when X = 19 AND Y = 41 else
"000000000000" when X = 20 AND Y = 41 else
"000000000000" when X = 21 AND Y = 41 else
"000000000000" when X = 22 AND Y = 41 else
"000000000000" when X = 23 AND Y = 41 else
"000000000000" when X = 24 AND Y = 41 else
"000000000000" when X = 25 AND Y = 41 else
"000000000000" when X = 26 AND Y = 41 else
"000000000000" when X = 27 AND Y = 41 else
"000000000000" when X = 28 AND Y = 41 else
"000000000000" when X = 29 AND Y = 41 else
"000000000000" when X = 30 AND Y = 41 else
"000000000000" when X = 31 AND Y = 41 else
"000000000000" when X = 32 AND Y = 41 else
"000000000000" when X = 33 AND Y = 41 else
"000000000000" when X = 34 AND Y = 41 else
"000000000000" when X = 35 AND Y = 41 else
"000000000000" when X = 36 AND Y = 41 else
"000000000000" when X = 37 AND Y = 41 else
"000000000000" when X = 38 AND Y = 41 else
"000000000000" when X = 39 AND Y = 41 else
"100010011101" when X = 40 AND Y = 41 else
"100010011101" when X = 41 AND Y = 41 else
"100010011101" when X = 42 AND Y = 41 else
"100010011101" when X = 43 AND Y = 41 else
"100010011101" when X = 44 AND Y = 41 else
"100010011101" when X = 45 AND Y = 41 else
"100010011101" when X = 46 AND Y = 41 else
"100010011101" when X = 47 AND Y = 41 else
"100010011101" when X = 48 AND Y = 41 else
"100010011101" when X = 49 AND Y = 41 else
"110111011111" when X = 50 AND Y = 41 else
"110111011111" when X = 51 AND Y = 41 else
"110111011111" when X = 52 AND Y = 41 else
"110111011111" when X = 53 AND Y = 41 else
"110111011111" when X = 54 AND Y = 41 else
"110111011111" when X = 55 AND Y = 41 else
"110111011111" when X = 56 AND Y = 41 else
"110111011111" when X = 57 AND Y = 41 else
"110111011111" when X = 58 AND Y = 41 else
"110111011111" when X = 59 AND Y = 41 else
"111111111111" when X = 60 AND Y = 41 else
"111111111111" when X = 61 AND Y = 41 else
"111111111111" when X = 62 AND Y = 41 else
"111111111111" when X = 63 AND Y = 41 else
"111111111111" when X = 64 AND Y = 41 else
"111111111111" when X = 65 AND Y = 41 else
"111111111111" when X = 66 AND Y = 41 else
"111111111111" when X = 67 AND Y = 41 else
"111111111111" when X = 68 AND Y = 41 else
"111111111111" when X = 69 AND Y = 41 else
"111111111111" when X = 70 AND Y = 41 else
"111111111111" when X = 71 AND Y = 41 else
"111111111111" when X = 72 AND Y = 41 else
"111111111111" when X = 73 AND Y = 41 else
"111111111111" when X = 74 AND Y = 41 else
"111111111111" when X = 75 AND Y = 41 else
"111111111111" when X = 76 AND Y = 41 else
"111111111111" when X = 77 AND Y = 41 else
"111111111111" when X = 78 AND Y = 41 else
"111111111111" when X = 79 AND Y = 41 else
"111111111111" when X = 80 AND Y = 41 else
"111111111111" when X = 81 AND Y = 41 else
"111111111111" when X = 82 AND Y = 41 else
"111111111111" when X = 83 AND Y = 41 else
"111111111111" when X = 84 AND Y = 41 else
"111111111111" when X = 85 AND Y = 41 else
"111111111111" when X = 86 AND Y = 41 else
"111111111111" when X = 87 AND Y = 41 else
"111111111111" when X = 88 AND Y = 41 else
"111111111111" when X = 89 AND Y = 41 else
"111111111111" when X = 90 AND Y = 41 else
"111111111111" when X = 91 AND Y = 41 else
"111111111111" when X = 92 AND Y = 41 else
"111111111111" when X = 93 AND Y = 41 else
"111111111111" when X = 94 AND Y = 41 else
"111111111111" when X = 95 AND Y = 41 else
"111111111111" when X = 96 AND Y = 41 else
"111111111111" when X = 97 AND Y = 41 else
"111111111111" when X = 98 AND Y = 41 else
"111111111111" when X = 99 AND Y = 41 else
"111111111111" when X = 100 AND Y = 41 else
"111111111111" when X = 101 AND Y = 41 else
"111111111111" when X = 102 AND Y = 41 else
"111111111111" when X = 103 AND Y = 41 else
"111111111111" when X = 104 AND Y = 41 else
"111111111111" when X = 105 AND Y = 41 else
"111111111111" when X = 106 AND Y = 41 else
"111111111111" when X = 107 AND Y = 41 else
"111111111111" when X = 108 AND Y = 41 else
"111111111111" when X = 109 AND Y = 41 else
"111111111111" when X = 110 AND Y = 41 else
"111111111111" when X = 111 AND Y = 41 else
"111111111111" when X = 112 AND Y = 41 else
"111111111111" when X = 113 AND Y = 41 else
"111111111111" when X = 114 AND Y = 41 else
"111111111111" when X = 115 AND Y = 41 else
"111111111111" when X = 116 AND Y = 41 else
"111111111111" when X = 117 AND Y = 41 else
"111111111111" when X = 118 AND Y = 41 else
"111111111111" when X = 119 AND Y = 41 else
"111111111111" when X = 120 AND Y = 41 else
"111111111111" when X = 121 AND Y = 41 else
"111111111111" when X = 122 AND Y = 41 else
"111111111111" when X = 123 AND Y = 41 else
"111111111111" when X = 124 AND Y = 41 else
"111111111111" when X = 125 AND Y = 41 else
"111111111111" when X = 126 AND Y = 41 else
"111111111111" when X = 127 AND Y = 41 else
"111111111111" when X = 128 AND Y = 41 else
"111111111111" when X = 129 AND Y = 41 else
"111111111111" when X = 130 AND Y = 41 else
"111111111111" when X = 131 AND Y = 41 else
"111111111111" when X = 132 AND Y = 41 else
"111111111111" when X = 133 AND Y = 41 else
"111111111111" when X = 134 AND Y = 41 else
"111111111111" when X = 135 AND Y = 41 else
"111111111111" when X = 136 AND Y = 41 else
"111111111111" when X = 137 AND Y = 41 else
"111111111111" when X = 138 AND Y = 41 else
"111111111111" when X = 139 AND Y = 41 else
"111111111111" when X = 140 AND Y = 41 else
"111111111111" when X = 141 AND Y = 41 else
"111111111111" when X = 142 AND Y = 41 else
"111111111111" when X = 143 AND Y = 41 else
"111111111111" when X = 144 AND Y = 41 else
"111111111111" when X = 145 AND Y = 41 else
"111111111111" when X = 146 AND Y = 41 else
"111111111111" when X = 147 AND Y = 41 else
"111111111111" when X = 148 AND Y = 41 else
"111111111111" when X = 149 AND Y = 41 else
"111111111111" when X = 150 AND Y = 41 else
"111111111111" when X = 151 AND Y = 41 else
"111111111111" when X = 152 AND Y = 41 else
"111111111111" when X = 153 AND Y = 41 else
"111111111111" when X = 154 AND Y = 41 else
"111111111111" when X = 155 AND Y = 41 else
"111111111111" when X = 156 AND Y = 41 else
"111111111111" when X = 157 AND Y = 41 else
"111111111111" when X = 158 AND Y = 41 else
"111111111111" when X = 159 AND Y = 41 else
"111111111111" when X = 160 AND Y = 41 else
"111111111111" when X = 161 AND Y = 41 else
"111111111111" when X = 162 AND Y = 41 else
"111111111111" when X = 163 AND Y = 41 else
"111111111111" when X = 164 AND Y = 41 else
"111111111111" when X = 165 AND Y = 41 else
"111111111111" when X = 166 AND Y = 41 else
"111111111111" when X = 167 AND Y = 41 else
"111111111111" when X = 168 AND Y = 41 else
"111111111111" when X = 169 AND Y = 41 else
"111111111111" when X = 170 AND Y = 41 else
"111111111111" when X = 171 AND Y = 41 else
"111111111111" when X = 172 AND Y = 41 else
"111111111111" when X = 173 AND Y = 41 else
"111111111111" when X = 174 AND Y = 41 else
"111111111111" when X = 175 AND Y = 41 else
"111111111111" when X = 176 AND Y = 41 else
"111111111111" when X = 177 AND Y = 41 else
"111111111111" when X = 178 AND Y = 41 else
"111111111111" when X = 179 AND Y = 41 else
"111111111111" when X = 180 AND Y = 41 else
"111111111111" when X = 181 AND Y = 41 else
"111111111111" when X = 182 AND Y = 41 else
"111111111111" when X = 183 AND Y = 41 else
"111111111111" when X = 184 AND Y = 41 else
"111111111111" when X = 185 AND Y = 41 else
"111111111111" when X = 186 AND Y = 41 else
"111111111111" when X = 187 AND Y = 41 else
"111111111111" when X = 188 AND Y = 41 else
"111111111111" when X = 189 AND Y = 41 else
"111111111111" when X = 190 AND Y = 41 else
"111111111111" when X = 191 AND Y = 41 else
"111111111111" when X = 192 AND Y = 41 else
"111111111111" when X = 193 AND Y = 41 else
"111111111111" when X = 194 AND Y = 41 else
"111111111111" when X = 195 AND Y = 41 else
"111111111111" when X = 196 AND Y = 41 else
"111111111111" when X = 197 AND Y = 41 else
"111111111111" when X = 198 AND Y = 41 else
"111111111111" when X = 199 AND Y = 41 else
"111111111111" when X = 200 AND Y = 41 else
"111111111111" when X = 201 AND Y = 41 else
"111111111111" when X = 202 AND Y = 41 else
"111111111111" when X = 203 AND Y = 41 else
"111111111111" when X = 204 AND Y = 41 else
"111111111111" when X = 205 AND Y = 41 else
"111111111111" when X = 206 AND Y = 41 else
"111111111111" when X = 207 AND Y = 41 else
"111111111111" when X = 208 AND Y = 41 else
"111111111111" when X = 209 AND Y = 41 else
"111111111111" when X = 210 AND Y = 41 else
"111111111111" when X = 211 AND Y = 41 else
"111111111111" when X = 212 AND Y = 41 else
"111111111111" when X = 213 AND Y = 41 else
"111111111111" when X = 214 AND Y = 41 else
"111111111111" when X = 215 AND Y = 41 else
"111111111111" when X = 216 AND Y = 41 else
"111111111111" when X = 217 AND Y = 41 else
"111111111111" when X = 218 AND Y = 41 else
"111111111111" when X = 219 AND Y = 41 else
"111111111111" when X = 220 AND Y = 41 else
"111111111111" when X = 221 AND Y = 41 else
"111111111111" when X = 222 AND Y = 41 else
"111111111111" when X = 223 AND Y = 41 else
"111111111111" when X = 224 AND Y = 41 else
"111111111111" when X = 225 AND Y = 41 else
"111111111111" when X = 226 AND Y = 41 else
"111111111111" when X = 227 AND Y = 41 else
"111111111111" when X = 228 AND Y = 41 else
"111111111111" when X = 229 AND Y = 41 else
"111111111111" when X = 230 AND Y = 41 else
"111111111111" when X = 231 AND Y = 41 else
"111111111111" when X = 232 AND Y = 41 else
"111111111111" when X = 233 AND Y = 41 else
"111111111111" when X = 234 AND Y = 41 else
"111111111111" when X = 235 AND Y = 41 else
"111111111111" when X = 236 AND Y = 41 else
"111111111111" when X = 237 AND Y = 41 else
"111111111111" when X = 238 AND Y = 41 else
"111111111111" when X = 239 AND Y = 41 else
"111111111111" when X = 240 AND Y = 41 else
"111111111111" when X = 241 AND Y = 41 else
"111111111111" when X = 242 AND Y = 41 else
"111111111111" when X = 243 AND Y = 41 else
"111111111111" when X = 244 AND Y = 41 else
"111111111111" when X = 245 AND Y = 41 else
"111111111111" when X = 246 AND Y = 41 else
"111111111111" when X = 247 AND Y = 41 else
"111111111111" when X = 248 AND Y = 41 else
"111111111111" when X = 249 AND Y = 41 else
"111111111111" when X = 250 AND Y = 41 else
"111111111111" when X = 251 AND Y = 41 else
"111111111111" when X = 252 AND Y = 41 else
"111111111111" when X = 253 AND Y = 41 else
"111111111111" when X = 254 AND Y = 41 else
"111111111111" when X = 255 AND Y = 41 else
"111111111111" when X = 256 AND Y = 41 else
"111111111111" when X = 257 AND Y = 41 else
"111111111111" when X = 258 AND Y = 41 else
"111111111111" when X = 259 AND Y = 41 else
"111111111111" when X = 260 AND Y = 41 else
"111111111111" when X = 261 AND Y = 41 else
"111111111111" when X = 262 AND Y = 41 else
"111111111111" when X = 263 AND Y = 41 else
"111111111111" when X = 264 AND Y = 41 else
"110111011111" when X = 265 AND Y = 41 else
"110111011111" when X = 266 AND Y = 41 else
"110111011111" when X = 267 AND Y = 41 else
"110111011111" when X = 268 AND Y = 41 else
"110111011111" when X = 269 AND Y = 41 else
"110111011111" when X = 270 AND Y = 41 else
"110111011111" when X = 271 AND Y = 41 else
"110111011111" when X = 272 AND Y = 41 else
"110111011111" when X = 273 AND Y = 41 else
"110111011111" when X = 274 AND Y = 41 else
"110111011111" when X = 275 AND Y = 41 else
"110111011111" when X = 276 AND Y = 41 else
"110111011111" when X = 277 AND Y = 41 else
"110111011111" when X = 278 AND Y = 41 else
"110111011111" when X = 279 AND Y = 41 else
"000000000000" when X = 280 AND Y = 41 else
"000000000000" when X = 281 AND Y = 41 else
"000000000000" when X = 282 AND Y = 41 else
"000000000000" when X = 283 AND Y = 41 else
"000000000000" when X = 284 AND Y = 41 else
"000000000000" when X = 285 AND Y = 41 else
"000000000000" when X = 286 AND Y = 41 else
"000000000000" when X = 287 AND Y = 41 else
"000000000000" when X = 288 AND Y = 41 else
"000000000000" when X = 289 AND Y = 41 else
"000000000000" when X = 290 AND Y = 41 else
"000000000000" when X = 291 AND Y = 41 else
"000000000000" when X = 292 AND Y = 41 else
"000000000000" when X = 293 AND Y = 41 else
"000000000000" when X = 294 AND Y = 41 else
"000000000000" when X = 295 AND Y = 41 else
"000000000000" when X = 296 AND Y = 41 else
"000000000000" when X = 297 AND Y = 41 else
"000000000000" when X = 298 AND Y = 41 else
"000000000000" when X = 299 AND Y = 41 else
"000000000000" when X = 300 AND Y = 41 else
"000000000000" when X = 301 AND Y = 41 else
"000000000000" when X = 302 AND Y = 41 else
"000000000000" when X = 303 AND Y = 41 else
"000000000000" when X = 304 AND Y = 41 else
"000000000000" when X = 305 AND Y = 41 else
"000000000000" when X = 306 AND Y = 41 else
"000000000000" when X = 307 AND Y = 41 else
"000000000000" when X = 308 AND Y = 41 else
"000000000000" when X = 309 AND Y = 41 else
"000000000000" when X = 310 AND Y = 41 else
"000000000000" when X = 311 AND Y = 41 else
"000000000000" when X = 312 AND Y = 41 else
"000000000000" when X = 313 AND Y = 41 else
"000000000000" when X = 314 AND Y = 41 else
"000000000000" when X = 315 AND Y = 41 else
"000000000000" when X = 316 AND Y = 41 else
"000000000000" when X = 317 AND Y = 41 else
"000000000000" when X = 318 AND Y = 41 else
"000000000000" when X = 319 AND Y = 41 else
"000000000000" when X = 320 AND Y = 41 else
"000000000000" when X = 321 AND Y = 41 else
"000000000000" when X = 322 AND Y = 41 else
"000000000000" when X = 323 AND Y = 41 else
"000000000000" when X = 324 AND Y = 41 else
"000000000000" when X = 0 AND Y = 42 else
"000000000000" when X = 1 AND Y = 42 else
"000000000000" when X = 2 AND Y = 42 else
"000000000000" when X = 3 AND Y = 42 else
"000000000000" when X = 4 AND Y = 42 else
"000000000000" when X = 5 AND Y = 42 else
"000000000000" when X = 6 AND Y = 42 else
"000000000000" when X = 7 AND Y = 42 else
"000000000000" when X = 8 AND Y = 42 else
"000000000000" when X = 9 AND Y = 42 else
"000000000000" when X = 10 AND Y = 42 else
"000000000000" when X = 11 AND Y = 42 else
"000000000000" when X = 12 AND Y = 42 else
"000000000000" when X = 13 AND Y = 42 else
"000000000000" when X = 14 AND Y = 42 else
"000000000000" when X = 15 AND Y = 42 else
"000000000000" when X = 16 AND Y = 42 else
"000000000000" when X = 17 AND Y = 42 else
"000000000000" when X = 18 AND Y = 42 else
"000000000000" when X = 19 AND Y = 42 else
"000000000000" when X = 20 AND Y = 42 else
"000000000000" when X = 21 AND Y = 42 else
"000000000000" when X = 22 AND Y = 42 else
"000000000000" when X = 23 AND Y = 42 else
"000000000000" when X = 24 AND Y = 42 else
"000000000000" when X = 25 AND Y = 42 else
"000000000000" when X = 26 AND Y = 42 else
"000000000000" when X = 27 AND Y = 42 else
"000000000000" when X = 28 AND Y = 42 else
"000000000000" when X = 29 AND Y = 42 else
"000000000000" when X = 30 AND Y = 42 else
"000000000000" when X = 31 AND Y = 42 else
"000000000000" when X = 32 AND Y = 42 else
"000000000000" when X = 33 AND Y = 42 else
"000000000000" when X = 34 AND Y = 42 else
"000000000000" when X = 35 AND Y = 42 else
"000000000000" when X = 36 AND Y = 42 else
"000000000000" when X = 37 AND Y = 42 else
"000000000000" when X = 38 AND Y = 42 else
"000000000000" when X = 39 AND Y = 42 else
"100010011101" when X = 40 AND Y = 42 else
"100010011101" when X = 41 AND Y = 42 else
"100010011101" when X = 42 AND Y = 42 else
"100010011101" when X = 43 AND Y = 42 else
"100010011101" when X = 44 AND Y = 42 else
"100010011101" when X = 45 AND Y = 42 else
"100010011101" when X = 46 AND Y = 42 else
"100010011101" when X = 47 AND Y = 42 else
"100010011101" when X = 48 AND Y = 42 else
"100010011101" when X = 49 AND Y = 42 else
"110111011111" when X = 50 AND Y = 42 else
"110111011111" when X = 51 AND Y = 42 else
"110111011111" when X = 52 AND Y = 42 else
"110111011111" when X = 53 AND Y = 42 else
"110111011111" when X = 54 AND Y = 42 else
"110111011111" when X = 55 AND Y = 42 else
"110111011111" when X = 56 AND Y = 42 else
"110111011111" when X = 57 AND Y = 42 else
"110111011111" when X = 58 AND Y = 42 else
"110111011111" when X = 59 AND Y = 42 else
"111111111111" when X = 60 AND Y = 42 else
"111111111111" when X = 61 AND Y = 42 else
"111111111111" when X = 62 AND Y = 42 else
"111111111111" when X = 63 AND Y = 42 else
"111111111111" when X = 64 AND Y = 42 else
"111111111111" when X = 65 AND Y = 42 else
"111111111111" when X = 66 AND Y = 42 else
"111111111111" when X = 67 AND Y = 42 else
"111111111111" when X = 68 AND Y = 42 else
"111111111111" when X = 69 AND Y = 42 else
"111111111111" when X = 70 AND Y = 42 else
"111111111111" when X = 71 AND Y = 42 else
"111111111111" when X = 72 AND Y = 42 else
"111111111111" when X = 73 AND Y = 42 else
"111111111111" when X = 74 AND Y = 42 else
"111111111111" when X = 75 AND Y = 42 else
"111111111111" when X = 76 AND Y = 42 else
"111111111111" when X = 77 AND Y = 42 else
"111111111111" when X = 78 AND Y = 42 else
"111111111111" when X = 79 AND Y = 42 else
"111111111111" when X = 80 AND Y = 42 else
"111111111111" when X = 81 AND Y = 42 else
"111111111111" when X = 82 AND Y = 42 else
"111111111111" when X = 83 AND Y = 42 else
"111111111111" when X = 84 AND Y = 42 else
"111111111111" when X = 85 AND Y = 42 else
"111111111111" when X = 86 AND Y = 42 else
"111111111111" when X = 87 AND Y = 42 else
"111111111111" when X = 88 AND Y = 42 else
"111111111111" when X = 89 AND Y = 42 else
"111111111111" when X = 90 AND Y = 42 else
"111111111111" when X = 91 AND Y = 42 else
"111111111111" when X = 92 AND Y = 42 else
"111111111111" when X = 93 AND Y = 42 else
"111111111111" when X = 94 AND Y = 42 else
"111111111111" when X = 95 AND Y = 42 else
"111111111111" when X = 96 AND Y = 42 else
"111111111111" when X = 97 AND Y = 42 else
"111111111111" when X = 98 AND Y = 42 else
"111111111111" when X = 99 AND Y = 42 else
"111111111111" when X = 100 AND Y = 42 else
"111111111111" when X = 101 AND Y = 42 else
"111111111111" when X = 102 AND Y = 42 else
"111111111111" when X = 103 AND Y = 42 else
"111111111111" when X = 104 AND Y = 42 else
"111111111111" when X = 105 AND Y = 42 else
"111111111111" when X = 106 AND Y = 42 else
"111111111111" when X = 107 AND Y = 42 else
"111111111111" when X = 108 AND Y = 42 else
"111111111111" when X = 109 AND Y = 42 else
"111111111111" when X = 110 AND Y = 42 else
"111111111111" when X = 111 AND Y = 42 else
"111111111111" when X = 112 AND Y = 42 else
"111111111111" when X = 113 AND Y = 42 else
"111111111111" when X = 114 AND Y = 42 else
"111111111111" when X = 115 AND Y = 42 else
"111111111111" when X = 116 AND Y = 42 else
"111111111111" when X = 117 AND Y = 42 else
"111111111111" when X = 118 AND Y = 42 else
"111111111111" when X = 119 AND Y = 42 else
"111111111111" when X = 120 AND Y = 42 else
"111111111111" when X = 121 AND Y = 42 else
"111111111111" when X = 122 AND Y = 42 else
"111111111111" when X = 123 AND Y = 42 else
"111111111111" when X = 124 AND Y = 42 else
"111111111111" when X = 125 AND Y = 42 else
"111111111111" when X = 126 AND Y = 42 else
"111111111111" when X = 127 AND Y = 42 else
"111111111111" when X = 128 AND Y = 42 else
"111111111111" when X = 129 AND Y = 42 else
"111111111111" when X = 130 AND Y = 42 else
"111111111111" when X = 131 AND Y = 42 else
"111111111111" when X = 132 AND Y = 42 else
"111111111111" when X = 133 AND Y = 42 else
"111111111111" when X = 134 AND Y = 42 else
"111111111111" when X = 135 AND Y = 42 else
"111111111111" when X = 136 AND Y = 42 else
"111111111111" when X = 137 AND Y = 42 else
"111111111111" when X = 138 AND Y = 42 else
"111111111111" when X = 139 AND Y = 42 else
"111111111111" when X = 140 AND Y = 42 else
"111111111111" when X = 141 AND Y = 42 else
"111111111111" when X = 142 AND Y = 42 else
"111111111111" when X = 143 AND Y = 42 else
"111111111111" when X = 144 AND Y = 42 else
"111111111111" when X = 145 AND Y = 42 else
"111111111111" when X = 146 AND Y = 42 else
"111111111111" when X = 147 AND Y = 42 else
"111111111111" when X = 148 AND Y = 42 else
"111111111111" when X = 149 AND Y = 42 else
"111111111111" when X = 150 AND Y = 42 else
"111111111111" when X = 151 AND Y = 42 else
"111111111111" when X = 152 AND Y = 42 else
"111111111111" when X = 153 AND Y = 42 else
"111111111111" when X = 154 AND Y = 42 else
"111111111111" when X = 155 AND Y = 42 else
"111111111111" when X = 156 AND Y = 42 else
"111111111111" when X = 157 AND Y = 42 else
"111111111111" when X = 158 AND Y = 42 else
"111111111111" when X = 159 AND Y = 42 else
"111111111111" when X = 160 AND Y = 42 else
"111111111111" when X = 161 AND Y = 42 else
"111111111111" when X = 162 AND Y = 42 else
"111111111111" when X = 163 AND Y = 42 else
"111111111111" when X = 164 AND Y = 42 else
"111111111111" when X = 165 AND Y = 42 else
"111111111111" when X = 166 AND Y = 42 else
"111111111111" when X = 167 AND Y = 42 else
"111111111111" when X = 168 AND Y = 42 else
"111111111111" when X = 169 AND Y = 42 else
"111111111111" when X = 170 AND Y = 42 else
"111111111111" when X = 171 AND Y = 42 else
"111111111111" when X = 172 AND Y = 42 else
"111111111111" when X = 173 AND Y = 42 else
"111111111111" when X = 174 AND Y = 42 else
"111111111111" when X = 175 AND Y = 42 else
"111111111111" when X = 176 AND Y = 42 else
"111111111111" when X = 177 AND Y = 42 else
"111111111111" when X = 178 AND Y = 42 else
"111111111111" when X = 179 AND Y = 42 else
"111111111111" when X = 180 AND Y = 42 else
"111111111111" when X = 181 AND Y = 42 else
"111111111111" when X = 182 AND Y = 42 else
"111111111111" when X = 183 AND Y = 42 else
"111111111111" when X = 184 AND Y = 42 else
"111111111111" when X = 185 AND Y = 42 else
"111111111111" when X = 186 AND Y = 42 else
"111111111111" when X = 187 AND Y = 42 else
"111111111111" when X = 188 AND Y = 42 else
"111111111111" when X = 189 AND Y = 42 else
"111111111111" when X = 190 AND Y = 42 else
"111111111111" when X = 191 AND Y = 42 else
"111111111111" when X = 192 AND Y = 42 else
"111111111111" when X = 193 AND Y = 42 else
"111111111111" when X = 194 AND Y = 42 else
"111111111111" when X = 195 AND Y = 42 else
"111111111111" when X = 196 AND Y = 42 else
"111111111111" when X = 197 AND Y = 42 else
"111111111111" when X = 198 AND Y = 42 else
"111111111111" when X = 199 AND Y = 42 else
"111111111111" when X = 200 AND Y = 42 else
"111111111111" when X = 201 AND Y = 42 else
"111111111111" when X = 202 AND Y = 42 else
"111111111111" when X = 203 AND Y = 42 else
"111111111111" when X = 204 AND Y = 42 else
"111111111111" when X = 205 AND Y = 42 else
"111111111111" when X = 206 AND Y = 42 else
"111111111111" when X = 207 AND Y = 42 else
"111111111111" when X = 208 AND Y = 42 else
"111111111111" when X = 209 AND Y = 42 else
"111111111111" when X = 210 AND Y = 42 else
"111111111111" when X = 211 AND Y = 42 else
"111111111111" when X = 212 AND Y = 42 else
"111111111111" when X = 213 AND Y = 42 else
"111111111111" when X = 214 AND Y = 42 else
"111111111111" when X = 215 AND Y = 42 else
"111111111111" when X = 216 AND Y = 42 else
"111111111111" when X = 217 AND Y = 42 else
"111111111111" when X = 218 AND Y = 42 else
"111111111111" when X = 219 AND Y = 42 else
"111111111111" when X = 220 AND Y = 42 else
"111111111111" when X = 221 AND Y = 42 else
"111111111111" when X = 222 AND Y = 42 else
"111111111111" when X = 223 AND Y = 42 else
"111111111111" when X = 224 AND Y = 42 else
"111111111111" when X = 225 AND Y = 42 else
"111111111111" when X = 226 AND Y = 42 else
"111111111111" when X = 227 AND Y = 42 else
"111111111111" when X = 228 AND Y = 42 else
"111111111111" when X = 229 AND Y = 42 else
"111111111111" when X = 230 AND Y = 42 else
"111111111111" when X = 231 AND Y = 42 else
"111111111111" when X = 232 AND Y = 42 else
"111111111111" when X = 233 AND Y = 42 else
"111111111111" when X = 234 AND Y = 42 else
"111111111111" when X = 235 AND Y = 42 else
"111111111111" when X = 236 AND Y = 42 else
"111111111111" when X = 237 AND Y = 42 else
"111111111111" when X = 238 AND Y = 42 else
"111111111111" when X = 239 AND Y = 42 else
"111111111111" when X = 240 AND Y = 42 else
"111111111111" when X = 241 AND Y = 42 else
"111111111111" when X = 242 AND Y = 42 else
"111111111111" when X = 243 AND Y = 42 else
"111111111111" when X = 244 AND Y = 42 else
"111111111111" when X = 245 AND Y = 42 else
"111111111111" when X = 246 AND Y = 42 else
"111111111111" when X = 247 AND Y = 42 else
"111111111111" when X = 248 AND Y = 42 else
"111111111111" when X = 249 AND Y = 42 else
"111111111111" when X = 250 AND Y = 42 else
"111111111111" when X = 251 AND Y = 42 else
"111111111111" when X = 252 AND Y = 42 else
"111111111111" when X = 253 AND Y = 42 else
"111111111111" when X = 254 AND Y = 42 else
"111111111111" when X = 255 AND Y = 42 else
"111111111111" when X = 256 AND Y = 42 else
"111111111111" when X = 257 AND Y = 42 else
"111111111111" when X = 258 AND Y = 42 else
"111111111111" when X = 259 AND Y = 42 else
"111111111111" when X = 260 AND Y = 42 else
"111111111111" when X = 261 AND Y = 42 else
"111111111111" when X = 262 AND Y = 42 else
"111111111111" when X = 263 AND Y = 42 else
"111111111111" when X = 264 AND Y = 42 else
"110111011111" when X = 265 AND Y = 42 else
"110111011111" when X = 266 AND Y = 42 else
"110111011111" when X = 267 AND Y = 42 else
"110111011111" when X = 268 AND Y = 42 else
"110111011111" when X = 269 AND Y = 42 else
"110111011111" when X = 270 AND Y = 42 else
"110111011111" when X = 271 AND Y = 42 else
"110111011111" when X = 272 AND Y = 42 else
"110111011111" when X = 273 AND Y = 42 else
"110111011111" when X = 274 AND Y = 42 else
"110111011111" when X = 275 AND Y = 42 else
"110111011111" when X = 276 AND Y = 42 else
"110111011111" when X = 277 AND Y = 42 else
"110111011111" when X = 278 AND Y = 42 else
"110111011111" when X = 279 AND Y = 42 else
"000000000000" when X = 280 AND Y = 42 else
"000000000000" when X = 281 AND Y = 42 else
"000000000000" when X = 282 AND Y = 42 else
"000000000000" when X = 283 AND Y = 42 else
"000000000000" when X = 284 AND Y = 42 else
"000000000000" when X = 285 AND Y = 42 else
"000000000000" when X = 286 AND Y = 42 else
"000000000000" when X = 287 AND Y = 42 else
"000000000000" when X = 288 AND Y = 42 else
"000000000000" when X = 289 AND Y = 42 else
"000000000000" when X = 290 AND Y = 42 else
"000000000000" when X = 291 AND Y = 42 else
"000000000000" when X = 292 AND Y = 42 else
"000000000000" when X = 293 AND Y = 42 else
"000000000000" when X = 294 AND Y = 42 else
"000000000000" when X = 295 AND Y = 42 else
"000000000000" when X = 296 AND Y = 42 else
"000000000000" when X = 297 AND Y = 42 else
"000000000000" when X = 298 AND Y = 42 else
"000000000000" when X = 299 AND Y = 42 else
"000000000000" when X = 300 AND Y = 42 else
"000000000000" when X = 301 AND Y = 42 else
"000000000000" when X = 302 AND Y = 42 else
"000000000000" when X = 303 AND Y = 42 else
"000000000000" when X = 304 AND Y = 42 else
"000000000000" when X = 305 AND Y = 42 else
"000000000000" when X = 306 AND Y = 42 else
"000000000000" when X = 307 AND Y = 42 else
"000000000000" when X = 308 AND Y = 42 else
"000000000000" when X = 309 AND Y = 42 else
"000000000000" when X = 310 AND Y = 42 else
"000000000000" when X = 311 AND Y = 42 else
"000000000000" when X = 312 AND Y = 42 else
"000000000000" when X = 313 AND Y = 42 else
"000000000000" when X = 314 AND Y = 42 else
"000000000000" when X = 315 AND Y = 42 else
"000000000000" when X = 316 AND Y = 42 else
"000000000000" when X = 317 AND Y = 42 else
"000000000000" when X = 318 AND Y = 42 else
"000000000000" when X = 319 AND Y = 42 else
"000000000000" when X = 320 AND Y = 42 else
"000000000000" when X = 321 AND Y = 42 else
"000000000000" when X = 322 AND Y = 42 else
"000000000000" when X = 323 AND Y = 42 else
"000000000000" when X = 324 AND Y = 42 else
"000000000000" when X = 0 AND Y = 43 else
"000000000000" when X = 1 AND Y = 43 else
"000000000000" when X = 2 AND Y = 43 else
"000000000000" when X = 3 AND Y = 43 else
"000000000000" when X = 4 AND Y = 43 else
"000000000000" when X = 5 AND Y = 43 else
"000000000000" when X = 6 AND Y = 43 else
"000000000000" when X = 7 AND Y = 43 else
"000000000000" when X = 8 AND Y = 43 else
"000000000000" when X = 9 AND Y = 43 else
"000000000000" when X = 10 AND Y = 43 else
"000000000000" when X = 11 AND Y = 43 else
"000000000000" when X = 12 AND Y = 43 else
"000000000000" when X = 13 AND Y = 43 else
"000000000000" when X = 14 AND Y = 43 else
"000000000000" when X = 15 AND Y = 43 else
"000000000000" when X = 16 AND Y = 43 else
"000000000000" when X = 17 AND Y = 43 else
"000000000000" when X = 18 AND Y = 43 else
"000000000000" when X = 19 AND Y = 43 else
"000000000000" when X = 20 AND Y = 43 else
"000000000000" when X = 21 AND Y = 43 else
"000000000000" when X = 22 AND Y = 43 else
"000000000000" when X = 23 AND Y = 43 else
"000000000000" when X = 24 AND Y = 43 else
"000000000000" when X = 25 AND Y = 43 else
"000000000000" when X = 26 AND Y = 43 else
"000000000000" when X = 27 AND Y = 43 else
"000000000000" when X = 28 AND Y = 43 else
"000000000000" when X = 29 AND Y = 43 else
"000000000000" when X = 30 AND Y = 43 else
"000000000000" when X = 31 AND Y = 43 else
"000000000000" when X = 32 AND Y = 43 else
"000000000000" when X = 33 AND Y = 43 else
"000000000000" when X = 34 AND Y = 43 else
"000000000000" when X = 35 AND Y = 43 else
"000000000000" when X = 36 AND Y = 43 else
"000000000000" when X = 37 AND Y = 43 else
"000000000000" when X = 38 AND Y = 43 else
"000000000000" when X = 39 AND Y = 43 else
"100010011101" when X = 40 AND Y = 43 else
"100010011101" when X = 41 AND Y = 43 else
"100010011101" when X = 42 AND Y = 43 else
"100010011101" when X = 43 AND Y = 43 else
"100010011101" when X = 44 AND Y = 43 else
"100010011101" when X = 45 AND Y = 43 else
"100010011101" when X = 46 AND Y = 43 else
"100010011101" when X = 47 AND Y = 43 else
"100010011101" when X = 48 AND Y = 43 else
"100010011101" when X = 49 AND Y = 43 else
"110111011111" when X = 50 AND Y = 43 else
"110111011111" when X = 51 AND Y = 43 else
"110111011111" when X = 52 AND Y = 43 else
"110111011111" when X = 53 AND Y = 43 else
"110111011111" when X = 54 AND Y = 43 else
"110111011111" when X = 55 AND Y = 43 else
"110111011111" when X = 56 AND Y = 43 else
"110111011111" when X = 57 AND Y = 43 else
"110111011111" when X = 58 AND Y = 43 else
"110111011111" when X = 59 AND Y = 43 else
"111111111111" when X = 60 AND Y = 43 else
"111111111111" when X = 61 AND Y = 43 else
"111111111111" when X = 62 AND Y = 43 else
"111111111111" when X = 63 AND Y = 43 else
"111111111111" when X = 64 AND Y = 43 else
"111111111111" when X = 65 AND Y = 43 else
"111111111111" when X = 66 AND Y = 43 else
"111111111111" when X = 67 AND Y = 43 else
"111111111111" when X = 68 AND Y = 43 else
"111111111111" when X = 69 AND Y = 43 else
"111111111111" when X = 70 AND Y = 43 else
"111111111111" when X = 71 AND Y = 43 else
"111111111111" when X = 72 AND Y = 43 else
"111111111111" when X = 73 AND Y = 43 else
"111111111111" when X = 74 AND Y = 43 else
"111111111111" when X = 75 AND Y = 43 else
"111111111111" when X = 76 AND Y = 43 else
"111111111111" when X = 77 AND Y = 43 else
"111111111111" when X = 78 AND Y = 43 else
"111111111111" when X = 79 AND Y = 43 else
"111111111111" when X = 80 AND Y = 43 else
"111111111111" when X = 81 AND Y = 43 else
"111111111111" when X = 82 AND Y = 43 else
"111111111111" when X = 83 AND Y = 43 else
"111111111111" when X = 84 AND Y = 43 else
"111111111111" when X = 85 AND Y = 43 else
"111111111111" when X = 86 AND Y = 43 else
"111111111111" when X = 87 AND Y = 43 else
"111111111111" when X = 88 AND Y = 43 else
"111111111111" when X = 89 AND Y = 43 else
"111111111111" when X = 90 AND Y = 43 else
"111111111111" when X = 91 AND Y = 43 else
"111111111111" when X = 92 AND Y = 43 else
"111111111111" when X = 93 AND Y = 43 else
"111111111111" when X = 94 AND Y = 43 else
"111111111111" when X = 95 AND Y = 43 else
"111111111111" when X = 96 AND Y = 43 else
"111111111111" when X = 97 AND Y = 43 else
"111111111111" when X = 98 AND Y = 43 else
"111111111111" when X = 99 AND Y = 43 else
"111111111111" when X = 100 AND Y = 43 else
"111111111111" when X = 101 AND Y = 43 else
"111111111111" when X = 102 AND Y = 43 else
"111111111111" when X = 103 AND Y = 43 else
"111111111111" when X = 104 AND Y = 43 else
"111111111111" when X = 105 AND Y = 43 else
"111111111111" when X = 106 AND Y = 43 else
"111111111111" when X = 107 AND Y = 43 else
"111111111111" when X = 108 AND Y = 43 else
"111111111111" when X = 109 AND Y = 43 else
"111111111111" when X = 110 AND Y = 43 else
"111111111111" when X = 111 AND Y = 43 else
"111111111111" when X = 112 AND Y = 43 else
"111111111111" when X = 113 AND Y = 43 else
"111111111111" when X = 114 AND Y = 43 else
"111111111111" when X = 115 AND Y = 43 else
"111111111111" when X = 116 AND Y = 43 else
"111111111111" when X = 117 AND Y = 43 else
"111111111111" when X = 118 AND Y = 43 else
"111111111111" when X = 119 AND Y = 43 else
"111111111111" when X = 120 AND Y = 43 else
"111111111111" when X = 121 AND Y = 43 else
"111111111111" when X = 122 AND Y = 43 else
"111111111111" when X = 123 AND Y = 43 else
"111111111111" when X = 124 AND Y = 43 else
"111111111111" when X = 125 AND Y = 43 else
"111111111111" when X = 126 AND Y = 43 else
"111111111111" when X = 127 AND Y = 43 else
"111111111111" when X = 128 AND Y = 43 else
"111111111111" when X = 129 AND Y = 43 else
"111111111111" when X = 130 AND Y = 43 else
"111111111111" when X = 131 AND Y = 43 else
"111111111111" when X = 132 AND Y = 43 else
"111111111111" when X = 133 AND Y = 43 else
"111111111111" when X = 134 AND Y = 43 else
"111111111111" when X = 135 AND Y = 43 else
"111111111111" when X = 136 AND Y = 43 else
"111111111111" when X = 137 AND Y = 43 else
"111111111111" when X = 138 AND Y = 43 else
"111111111111" when X = 139 AND Y = 43 else
"111111111111" when X = 140 AND Y = 43 else
"111111111111" when X = 141 AND Y = 43 else
"111111111111" when X = 142 AND Y = 43 else
"111111111111" when X = 143 AND Y = 43 else
"111111111111" when X = 144 AND Y = 43 else
"111111111111" when X = 145 AND Y = 43 else
"111111111111" when X = 146 AND Y = 43 else
"111111111111" when X = 147 AND Y = 43 else
"111111111111" when X = 148 AND Y = 43 else
"111111111111" when X = 149 AND Y = 43 else
"111111111111" when X = 150 AND Y = 43 else
"111111111111" when X = 151 AND Y = 43 else
"111111111111" when X = 152 AND Y = 43 else
"111111111111" when X = 153 AND Y = 43 else
"111111111111" when X = 154 AND Y = 43 else
"111111111111" when X = 155 AND Y = 43 else
"111111111111" when X = 156 AND Y = 43 else
"111111111111" when X = 157 AND Y = 43 else
"111111111111" when X = 158 AND Y = 43 else
"111111111111" when X = 159 AND Y = 43 else
"111111111111" when X = 160 AND Y = 43 else
"111111111111" when X = 161 AND Y = 43 else
"111111111111" when X = 162 AND Y = 43 else
"111111111111" when X = 163 AND Y = 43 else
"111111111111" when X = 164 AND Y = 43 else
"111111111111" when X = 165 AND Y = 43 else
"111111111111" when X = 166 AND Y = 43 else
"111111111111" when X = 167 AND Y = 43 else
"111111111111" when X = 168 AND Y = 43 else
"111111111111" when X = 169 AND Y = 43 else
"111111111111" when X = 170 AND Y = 43 else
"111111111111" when X = 171 AND Y = 43 else
"111111111111" when X = 172 AND Y = 43 else
"111111111111" when X = 173 AND Y = 43 else
"111111111111" when X = 174 AND Y = 43 else
"111111111111" when X = 175 AND Y = 43 else
"111111111111" when X = 176 AND Y = 43 else
"111111111111" when X = 177 AND Y = 43 else
"111111111111" when X = 178 AND Y = 43 else
"111111111111" when X = 179 AND Y = 43 else
"111111111111" when X = 180 AND Y = 43 else
"111111111111" when X = 181 AND Y = 43 else
"111111111111" when X = 182 AND Y = 43 else
"111111111111" when X = 183 AND Y = 43 else
"111111111111" when X = 184 AND Y = 43 else
"111111111111" when X = 185 AND Y = 43 else
"111111111111" when X = 186 AND Y = 43 else
"111111111111" when X = 187 AND Y = 43 else
"111111111111" when X = 188 AND Y = 43 else
"111111111111" when X = 189 AND Y = 43 else
"111111111111" when X = 190 AND Y = 43 else
"111111111111" when X = 191 AND Y = 43 else
"111111111111" when X = 192 AND Y = 43 else
"111111111111" when X = 193 AND Y = 43 else
"111111111111" when X = 194 AND Y = 43 else
"111111111111" when X = 195 AND Y = 43 else
"111111111111" when X = 196 AND Y = 43 else
"111111111111" when X = 197 AND Y = 43 else
"111111111111" when X = 198 AND Y = 43 else
"111111111111" when X = 199 AND Y = 43 else
"111111111111" when X = 200 AND Y = 43 else
"111111111111" when X = 201 AND Y = 43 else
"111111111111" when X = 202 AND Y = 43 else
"111111111111" when X = 203 AND Y = 43 else
"111111111111" when X = 204 AND Y = 43 else
"111111111111" when X = 205 AND Y = 43 else
"111111111111" when X = 206 AND Y = 43 else
"111111111111" when X = 207 AND Y = 43 else
"111111111111" when X = 208 AND Y = 43 else
"111111111111" when X = 209 AND Y = 43 else
"111111111111" when X = 210 AND Y = 43 else
"111111111111" when X = 211 AND Y = 43 else
"111111111111" when X = 212 AND Y = 43 else
"111111111111" when X = 213 AND Y = 43 else
"111111111111" when X = 214 AND Y = 43 else
"111111111111" when X = 215 AND Y = 43 else
"111111111111" when X = 216 AND Y = 43 else
"111111111111" when X = 217 AND Y = 43 else
"111111111111" when X = 218 AND Y = 43 else
"111111111111" when X = 219 AND Y = 43 else
"111111111111" when X = 220 AND Y = 43 else
"111111111111" when X = 221 AND Y = 43 else
"111111111111" when X = 222 AND Y = 43 else
"111111111111" when X = 223 AND Y = 43 else
"111111111111" when X = 224 AND Y = 43 else
"111111111111" when X = 225 AND Y = 43 else
"111111111111" when X = 226 AND Y = 43 else
"111111111111" when X = 227 AND Y = 43 else
"111111111111" when X = 228 AND Y = 43 else
"111111111111" when X = 229 AND Y = 43 else
"111111111111" when X = 230 AND Y = 43 else
"111111111111" when X = 231 AND Y = 43 else
"111111111111" when X = 232 AND Y = 43 else
"111111111111" when X = 233 AND Y = 43 else
"111111111111" when X = 234 AND Y = 43 else
"111111111111" when X = 235 AND Y = 43 else
"111111111111" when X = 236 AND Y = 43 else
"111111111111" when X = 237 AND Y = 43 else
"111111111111" when X = 238 AND Y = 43 else
"111111111111" when X = 239 AND Y = 43 else
"111111111111" when X = 240 AND Y = 43 else
"111111111111" when X = 241 AND Y = 43 else
"111111111111" when X = 242 AND Y = 43 else
"111111111111" when X = 243 AND Y = 43 else
"111111111111" when X = 244 AND Y = 43 else
"111111111111" when X = 245 AND Y = 43 else
"111111111111" when X = 246 AND Y = 43 else
"111111111111" when X = 247 AND Y = 43 else
"111111111111" when X = 248 AND Y = 43 else
"111111111111" when X = 249 AND Y = 43 else
"111111111111" when X = 250 AND Y = 43 else
"111111111111" when X = 251 AND Y = 43 else
"111111111111" when X = 252 AND Y = 43 else
"111111111111" when X = 253 AND Y = 43 else
"111111111111" when X = 254 AND Y = 43 else
"111111111111" when X = 255 AND Y = 43 else
"111111111111" when X = 256 AND Y = 43 else
"111111111111" when X = 257 AND Y = 43 else
"111111111111" when X = 258 AND Y = 43 else
"111111111111" when X = 259 AND Y = 43 else
"111111111111" when X = 260 AND Y = 43 else
"111111111111" when X = 261 AND Y = 43 else
"111111111111" when X = 262 AND Y = 43 else
"111111111111" when X = 263 AND Y = 43 else
"111111111111" when X = 264 AND Y = 43 else
"110111011111" when X = 265 AND Y = 43 else
"110111011111" when X = 266 AND Y = 43 else
"110111011111" when X = 267 AND Y = 43 else
"110111011111" when X = 268 AND Y = 43 else
"110111011111" when X = 269 AND Y = 43 else
"110111011111" when X = 270 AND Y = 43 else
"110111011111" when X = 271 AND Y = 43 else
"110111011111" when X = 272 AND Y = 43 else
"110111011111" when X = 273 AND Y = 43 else
"110111011111" when X = 274 AND Y = 43 else
"110111011111" when X = 275 AND Y = 43 else
"110111011111" when X = 276 AND Y = 43 else
"110111011111" when X = 277 AND Y = 43 else
"110111011111" when X = 278 AND Y = 43 else
"110111011111" when X = 279 AND Y = 43 else
"000000000000" when X = 280 AND Y = 43 else
"000000000000" when X = 281 AND Y = 43 else
"000000000000" when X = 282 AND Y = 43 else
"000000000000" when X = 283 AND Y = 43 else
"000000000000" when X = 284 AND Y = 43 else
"000000000000" when X = 285 AND Y = 43 else
"000000000000" when X = 286 AND Y = 43 else
"000000000000" when X = 287 AND Y = 43 else
"000000000000" when X = 288 AND Y = 43 else
"000000000000" when X = 289 AND Y = 43 else
"000000000000" when X = 290 AND Y = 43 else
"000000000000" when X = 291 AND Y = 43 else
"000000000000" when X = 292 AND Y = 43 else
"000000000000" when X = 293 AND Y = 43 else
"000000000000" when X = 294 AND Y = 43 else
"000000000000" when X = 295 AND Y = 43 else
"000000000000" when X = 296 AND Y = 43 else
"000000000000" when X = 297 AND Y = 43 else
"000000000000" when X = 298 AND Y = 43 else
"000000000000" when X = 299 AND Y = 43 else
"000000000000" when X = 300 AND Y = 43 else
"000000000000" when X = 301 AND Y = 43 else
"000000000000" when X = 302 AND Y = 43 else
"000000000000" when X = 303 AND Y = 43 else
"000000000000" when X = 304 AND Y = 43 else
"000000000000" when X = 305 AND Y = 43 else
"000000000000" when X = 306 AND Y = 43 else
"000000000000" when X = 307 AND Y = 43 else
"000000000000" when X = 308 AND Y = 43 else
"000000000000" when X = 309 AND Y = 43 else
"000000000000" when X = 310 AND Y = 43 else
"000000000000" when X = 311 AND Y = 43 else
"000000000000" when X = 312 AND Y = 43 else
"000000000000" when X = 313 AND Y = 43 else
"000000000000" when X = 314 AND Y = 43 else
"000000000000" when X = 315 AND Y = 43 else
"000000000000" when X = 316 AND Y = 43 else
"000000000000" when X = 317 AND Y = 43 else
"000000000000" when X = 318 AND Y = 43 else
"000000000000" when X = 319 AND Y = 43 else
"000000000000" when X = 320 AND Y = 43 else
"000000000000" when X = 321 AND Y = 43 else
"000000000000" when X = 322 AND Y = 43 else
"000000000000" when X = 323 AND Y = 43 else
"000000000000" when X = 324 AND Y = 43 else
"000000000000" when X = 0 AND Y = 44 else
"000000000000" when X = 1 AND Y = 44 else
"000000000000" when X = 2 AND Y = 44 else
"000000000000" when X = 3 AND Y = 44 else
"000000000000" when X = 4 AND Y = 44 else
"000000000000" when X = 5 AND Y = 44 else
"000000000000" when X = 6 AND Y = 44 else
"000000000000" when X = 7 AND Y = 44 else
"000000000000" when X = 8 AND Y = 44 else
"000000000000" when X = 9 AND Y = 44 else
"000000000000" when X = 10 AND Y = 44 else
"000000000000" when X = 11 AND Y = 44 else
"000000000000" when X = 12 AND Y = 44 else
"000000000000" when X = 13 AND Y = 44 else
"000000000000" when X = 14 AND Y = 44 else
"000000000000" when X = 15 AND Y = 44 else
"000000000000" when X = 16 AND Y = 44 else
"000000000000" when X = 17 AND Y = 44 else
"000000000000" when X = 18 AND Y = 44 else
"000000000000" when X = 19 AND Y = 44 else
"000000000000" when X = 20 AND Y = 44 else
"000000000000" when X = 21 AND Y = 44 else
"000000000000" when X = 22 AND Y = 44 else
"000000000000" when X = 23 AND Y = 44 else
"000000000000" when X = 24 AND Y = 44 else
"000000000000" when X = 25 AND Y = 44 else
"000000000000" when X = 26 AND Y = 44 else
"000000000000" when X = 27 AND Y = 44 else
"000000000000" when X = 28 AND Y = 44 else
"000000000000" when X = 29 AND Y = 44 else
"000000000000" when X = 30 AND Y = 44 else
"000000000000" when X = 31 AND Y = 44 else
"000000000000" when X = 32 AND Y = 44 else
"000000000000" when X = 33 AND Y = 44 else
"000000000000" when X = 34 AND Y = 44 else
"000000000000" when X = 35 AND Y = 44 else
"000000000000" when X = 36 AND Y = 44 else
"000000000000" when X = 37 AND Y = 44 else
"000000000000" when X = 38 AND Y = 44 else
"000000000000" when X = 39 AND Y = 44 else
"100010011101" when X = 40 AND Y = 44 else
"100010011101" when X = 41 AND Y = 44 else
"100010011101" when X = 42 AND Y = 44 else
"100010011101" when X = 43 AND Y = 44 else
"100010011101" when X = 44 AND Y = 44 else
"100010011101" when X = 45 AND Y = 44 else
"100010011101" when X = 46 AND Y = 44 else
"100010011101" when X = 47 AND Y = 44 else
"100010011101" when X = 48 AND Y = 44 else
"100010011101" when X = 49 AND Y = 44 else
"110111011111" when X = 50 AND Y = 44 else
"110111011111" when X = 51 AND Y = 44 else
"110111011111" when X = 52 AND Y = 44 else
"110111011111" when X = 53 AND Y = 44 else
"110111011111" when X = 54 AND Y = 44 else
"110111011111" when X = 55 AND Y = 44 else
"110111011111" when X = 56 AND Y = 44 else
"110111011111" when X = 57 AND Y = 44 else
"110111011111" when X = 58 AND Y = 44 else
"110111011111" when X = 59 AND Y = 44 else
"111111111111" when X = 60 AND Y = 44 else
"111111111111" when X = 61 AND Y = 44 else
"111111111111" when X = 62 AND Y = 44 else
"111111111111" when X = 63 AND Y = 44 else
"111111111111" when X = 64 AND Y = 44 else
"111111111111" when X = 65 AND Y = 44 else
"111111111111" when X = 66 AND Y = 44 else
"111111111111" when X = 67 AND Y = 44 else
"111111111111" when X = 68 AND Y = 44 else
"111111111111" when X = 69 AND Y = 44 else
"111111111111" when X = 70 AND Y = 44 else
"111111111111" when X = 71 AND Y = 44 else
"111111111111" when X = 72 AND Y = 44 else
"111111111111" when X = 73 AND Y = 44 else
"111111111111" when X = 74 AND Y = 44 else
"111111111111" when X = 75 AND Y = 44 else
"111111111111" when X = 76 AND Y = 44 else
"111111111111" when X = 77 AND Y = 44 else
"111111111111" when X = 78 AND Y = 44 else
"111111111111" when X = 79 AND Y = 44 else
"111111111111" when X = 80 AND Y = 44 else
"111111111111" when X = 81 AND Y = 44 else
"111111111111" when X = 82 AND Y = 44 else
"111111111111" when X = 83 AND Y = 44 else
"111111111111" when X = 84 AND Y = 44 else
"111111111111" when X = 85 AND Y = 44 else
"111111111111" when X = 86 AND Y = 44 else
"111111111111" when X = 87 AND Y = 44 else
"111111111111" when X = 88 AND Y = 44 else
"111111111111" when X = 89 AND Y = 44 else
"111111111111" when X = 90 AND Y = 44 else
"111111111111" when X = 91 AND Y = 44 else
"111111111111" when X = 92 AND Y = 44 else
"111111111111" when X = 93 AND Y = 44 else
"111111111111" when X = 94 AND Y = 44 else
"111111111111" when X = 95 AND Y = 44 else
"111111111111" when X = 96 AND Y = 44 else
"111111111111" when X = 97 AND Y = 44 else
"111111111111" when X = 98 AND Y = 44 else
"111111111111" when X = 99 AND Y = 44 else
"111111111111" when X = 100 AND Y = 44 else
"111111111111" when X = 101 AND Y = 44 else
"111111111111" when X = 102 AND Y = 44 else
"111111111111" when X = 103 AND Y = 44 else
"111111111111" when X = 104 AND Y = 44 else
"111111111111" when X = 105 AND Y = 44 else
"111111111111" when X = 106 AND Y = 44 else
"111111111111" when X = 107 AND Y = 44 else
"111111111111" when X = 108 AND Y = 44 else
"111111111111" when X = 109 AND Y = 44 else
"111111111111" when X = 110 AND Y = 44 else
"111111111111" when X = 111 AND Y = 44 else
"111111111111" when X = 112 AND Y = 44 else
"111111111111" when X = 113 AND Y = 44 else
"111111111111" when X = 114 AND Y = 44 else
"111111111111" when X = 115 AND Y = 44 else
"111111111111" when X = 116 AND Y = 44 else
"111111111111" when X = 117 AND Y = 44 else
"111111111111" when X = 118 AND Y = 44 else
"111111111111" when X = 119 AND Y = 44 else
"111111111111" when X = 120 AND Y = 44 else
"111111111111" when X = 121 AND Y = 44 else
"111111111111" when X = 122 AND Y = 44 else
"111111111111" when X = 123 AND Y = 44 else
"111111111111" when X = 124 AND Y = 44 else
"111111111111" when X = 125 AND Y = 44 else
"111111111111" when X = 126 AND Y = 44 else
"111111111111" when X = 127 AND Y = 44 else
"111111111111" when X = 128 AND Y = 44 else
"111111111111" when X = 129 AND Y = 44 else
"111111111111" when X = 130 AND Y = 44 else
"111111111111" when X = 131 AND Y = 44 else
"111111111111" when X = 132 AND Y = 44 else
"111111111111" when X = 133 AND Y = 44 else
"111111111111" when X = 134 AND Y = 44 else
"111111111111" when X = 135 AND Y = 44 else
"111111111111" when X = 136 AND Y = 44 else
"111111111111" when X = 137 AND Y = 44 else
"111111111111" when X = 138 AND Y = 44 else
"111111111111" when X = 139 AND Y = 44 else
"111111111111" when X = 140 AND Y = 44 else
"111111111111" when X = 141 AND Y = 44 else
"111111111111" when X = 142 AND Y = 44 else
"111111111111" when X = 143 AND Y = 44 else
"111111111111" when X = 144 AND Y = 44 else
"111111111111" when X = 145 AND Y = 44 else
"111111111111" when X = 146 AND Y = 44 else
"111111111111" when X = 147 AND Y = 44 else
"111111111111" when X = 148 AND Y = 44 else
"111111111111" when X = 149 AND Y = 44 else
"111111111111" when X = 150 AND Y = 44 else
"111111111111" when X = 151 AND Y = 44 else
"111111111111" when X = 152 AND Y = 44 else
"111111111111" when X = 153 AND Y = 44 else
"111111111111" when X = 154 AND Y = 44 else
"111111111111" when X = 155 AND Y = 44 else
"111111111111" when X = 156 AND Y = 44 else
"111111111111" when X = 157 AND Y = 44 else
"111111111111" when X = 158 AND Y = 44 else
"111111111111" when X = 159 AND Y = 44 else
"111111111111" when X = 160 AND Y = 44 else
"111111111111" when X = 161 AND Y = 44 else
"111111111111" when X = 162 AND Y = 44 else
"111111111111" when X = 163 AND Y = 44 else
"111111111111" when X = 164 AND Y = 44 else
"111111111111" when X = 165 AND Y = 44 else
"111111111111" when X = 166 AND Y = 44 else
"111111111111" when X = 167 AND Y = 44 else
"111111111111" when X = 168 AND Y = 44 else
"111111111111" when X = 169 AND Y = 44 else
"111111111111" when X = 170 AND Y = 44 else
"111111111111" when X = 171 AND Y = 44 else
"111111111111" when X = 172 AND Y = 44 else
"111111111111" when X = 173 AND Y = 44 else
"111111111111" when X = 174 AND Y = 44 else
"111111111111" when X = 175 AND Y = 44 else
"111111111111" when X = 176 AND Y = 44 else
"111111111111" when X = 177 AND Y = 44 else
"111111111111" when X = 178 AND Y = 44 else
"111111111111" when X = 179 AND Y = 44 else
"111111111111" when X = 180 AND Y = 44 else
"111111111111" when X = 181 AND Y = 44 else
"111111111111" when X = 182 AND Y = 44 else
"111111111111" when X = 183 AND Y = 44 else
"111111111111" when X = 184 AND Y = 44 else
"111111111111" when X = 185 AND Y = 44 else
"111111111111" when X = 186 AND Y = 44 else
"111111111111" when X = 187 AND Y = 44 else
"111111111111" when X = 188 AND Y = 44 else
"111111111111" when X = 189 AND Y = 44 else
"111111111111" when X = 190 AND Y = 44 else
"111111111111" when X = 191 AND Y = 44 else
"111111111111" when X = 192 AND Y = 44 else
"111111111111" when X = 193 AND Y = 44 else
"111111111111" when X = 194 AND Y = 44 else
"111111111111" when X = 195 AND Y = 44 else
"111111111111" when X = 196 AND Y = 44 else
"111111111111" when X = 197 AND Y = 44 else
"111111111111" when X = 198 AND Y = 44 else
"111111111111" when X = 199 AND Y = 44 else
"111111111111" when X = 200 AND Y = 44 else
"111111111111" when X = 201 AND Y = 44 else
"111111111111" when X = 202 AND Y = 44 else
"111111111111" when X = 203 AND Y = 44 else
"111111111111" when X = 204 AND Y = 44 else
"111111111111" when X = 205 AND Y = 44 else
"111111111111" when X = 206 AND Y = 44 else
"111111111111" when X = 207 AND Y = 44 else
"111111111111" when X = 208 AND Y = 44 else
"111111111111" when X = 209 AND Y = 44 else
"111111111111" when X = 210 AND Y = 44 else
"111111111111" when X = 211 AND Y = 44 else
"111111111111" when X = 212 AND Y = 44 else
"111111111111" when X = 213 AND Y = 44 else
"111111111111" when X = 214 AND Y = 44 else
"111111111111" when X = 215 AND Y = 44 else
"111111111111" when X = 216 AND Y = 44 else
"111111111111" when X = 217 AND Y = 44 else
"111111111111" when X = 218 AND Y = 44 else
"111111111111" when X = 219 AND Y = 44 else
"111111111111" when X = 220 AND Y = 44 else
"111111111111" when X = 221 AND Y = 44 else
"111111111111" when X = 222 AND Y = 44 else
"111111111111" when X = 223 AND Y = 44 else
"111111111111" when X = 224 AND Y = 44 else
"111111111111" when X = 225 AND Y = 44 else
"111111111111" when X = 226 AND Y = 44 else
"111111111111" when X = 227 AND Y = 44 else
"111111111111" when X = 228 AND Y = 44 else
"111111111111" when X = 229 AND Y = 44 else
"111111111111" when X = 230 AND Y = 44 else
"111111111111" when X = 231 AND Y = 44 else
"111111111111" when X = 232 AND Y = 44 else
"111111111111" when X = 233 AND Y = 44 else
"111111111111" when X = 234 AND Y = 44 else
"111111111111" when X = 235 AND Y = 44 else
"111111111111" when X = 236 AND Y = 44 else
"111111111111" when X = 237 AND Y = 44 else
"111111111111" when X = 238 AND Y = 44 else
"111111111111" when X = 239 AND Y = 44 else
"111111111111" when X = 240 AND Y = 44 else
"111111111111" when X = 241 AND Y = 44 else
"111111111111" when X = 242 AND Y = 44 else
"111111111111" when X = 243 AND Y = 44 else
"111111111111" when X = 244 AND Y = 44 else
"111111111111" when X = 245 AND Y = 44 else
"111111111111" when X = 246 AND Y = 44 else
"111111111111" when X = 247 AND Y = 44 else
"111111111111" when X = 248 AND Y = 44 else
"111111111111" when X = 249 AND Y = 44 else
"111111111111" when X = 250 AND Y = 44 else
"111111111111" when X = 251 AND Y = 44 else
"111111111111" when X = 252 AND Y = 44 else
"111111111111" when X = 253 AND Y = 44 else
"111111111111" when X = 254 AND Y = 44 else
"111111111111" when X = 255 AND Y = 44 else
"111111111111" when X = 256 AND Y = 44 else
"111111111111" when X = 257 AND Y = 44 else
"111111111111" when X = 258 AND Y = 44 else
"111111111111" when X = 259 AND Y = 44 else
"111111111111" when X = 260 AND Y = 44 else
"111111111111" when X = 261 AND Y = 44 else
"111111111111" when X = 262 AND Y = 44 else
"111111111111" when X = 263 AND Y = 44 else
"111111111111" when X = 264 AND Y = 44 else
"110111011111" when X = 265 AND Y = 44 else
"110111011111" when X = 266 AND Y = 44 else
"110111011111" when X = 267 AND Y = 44 else
"110111011111" when X = 268 AND Y = 44 else
"110111011111" when X = 269 AND Y = 44 else
"110111011111" when X = 270 AND Y = 44 else
"110111011111" when X = 271 AND Y = 44 else
"110111011111" when X = 272 AND Y = 44 else
"110111011111" when X = 273 AND Y = 44 else
"110111011111" when X = 274 AND Y = 44 else
"110111011111" when X = 275 AND Y = 44 else
"110111011111" when X = 276 AND Y = 44 else
"110111011111" when X = 277 AND Y = 44 else
"110111011111" when X = 278 AND Y = 44 else
"110111011111" when X = 279 AND Y = 44 else
"000000000000" when X = 280 AND Y = 44 else
"000000000000" when X = 281 AND Y = 44 else
"000000000000" when X = 282 AND Y = 44 else
"000000000000" when X = 283 AND Y = 44 else
"000000000000" when X = 284 AND Y = 44 else
"000000000000" when X = 285 AND Y = 44 else
"000000000000" when X = 286 AND Y = 44 else
"000000000000" when X = 287 AND Y = 44 else
"000000000000" when X = 288 AND Y = 44 else
"000000000000" when X = 289 AND Y = 44 else
"000000000000" when X = 290 AND Y = 44 else
"000000000000" when X = 291 AND Y = 44 else
"000000000000" when X = 292 AND Y = 44 else
"000000000000" when X = 293 AND Y = 44 else
"000000000000" when X = 294 AND Y = 44 else
"000000000000" when X = 295 AND Y = 44 else
"000000000000" when X = 296 AND Y = 44 else
"000000000000" when X = 297 AND Y = 44 else
"000000000000" when X = 298 AND Y = 44 else
"000000000000" when X = 299 AND Y = 44 else
"000000000000" when X = 300 AND Y = 44 else
"000000000000" when X = 301 AND Y = 44 else
"000000000000" when X = 302 AND Y = 44 else
"000000000000" when X = 303 AND Y = 44 else
"000000000000" when X = 304 AND Y = 44 else
"000000000000" when X = 305 AND Y = 44 else
"000000000000" when X = 306 AND Y = 44 else
"000000000000" when X = 307 AND Y = 44 else
"000000000000" when X = 308 AND Y = 44 else
"000000000000" when X = 309 AND Y = 44 else
"000000000000" when X = 310 AND Y = 44 else
"000000000000" when X = 311 AND Y = 44 else
"000000000000" when X = 312 AND Y = 44 else
"000000000000" when X = 313 AND Y = 44 else
"000000000000" when X = 314 AND Y = 44 else
"000000000000" when X = 315 AND Y = 44 else
"000000000000" when X = 316 AND Y = 44 else
"000000000000" when X = 317 AND Y = 44 else
"000000000000" when X = 318 AND Y = 44 else
"000000000000" when X = 319 AND Y = 44 else
"000000000000" when X = 320 AND Y = 44 else
"000000000000" when X = 321 AND Y = 44 else
"000000000000" when X = 322 AND Y = 44 else
"000000000000" when X = 323 AND Y = 44 else
"000000000000" when X = 324 AND Y = 44 else
"000000000000" when X = 0 AND Y = 45 else
"000000000000" when X = 1 AND Y = 45 else
"000000000000" when X = 2 AND Y = 45 else
"000000000000" when X = 3 AND Y = 45 else
"000000000000" when X = 4 AND Y = 45 else
"000000000000" when X = 5 AND Y = 45 else
"000000000000" when X = 6 AND Y = 45 else
"000000000000" when X = 7 AND Y = 45 else
"000000000000" when X = 8 AND Y = 45 else
"000000000000" when X = 9 AND Y = 45 else
"000000000000" when X = 10 AND Y = 45 else
"000000000000" when X = 11 AND Y = 45 else
"000000000000" when X = 12 AND Y = 45 else
"000000000000" when X = 13 AND Y = 45 else
"000000000000" when X = 14 AND Y = 45 else
"000000000000" when X = 15 AND Y = 45 else
"000000000000" when X = 16 AND Y = 45 else
"000000000000" when X = 17 AND Y = 45 else
"000000000000" when X = 18 AND Y = 45 else
"000000000000" when X = 19 AND Y = 45 else
"000000000000" when X = 20 AND Y = 45 else
"000000000000" when X = 21 AND Y = 45 else
"000000000000" when X = 22 AND Y = 45 else
"000000000000" when X = 23 AND Y = 45 else
"000000000000" when X = 24 AND Y = 45 else
"000000000000" when X = 25 AND Y = 45 else
"000000000000" when X = 26 AND Y = 45 else
"000000000000" when X = 27 AND Y = 45 else
"000000000000" when X = 28 AND Y = 45 else
"000000000000" when X = 29 AND Y = 45 else
"000000000000" when X = 30 AND Y = 45 else
"000000000000" when X = 31 AND Y = 45 else
"000000000000" when X = 32 AND Y = 45 else
"000000000000" when X = 33 AND Y = 45 else
"000000000000" when X = 34 AND Y = 45 else
"000000000000" when X = 35 AND Y = 45 else
"000000000000" when X = 36 AND Y = 45 else
"000000000000" when X = 37 AND Y = 45 else
"000000000000" when X = 38 AND Y = 45 else
"000000000000" when X = 39 AND Y = 45 else
"100010011101" when X = 40 AND Y = 45 else
"100010011101" when X = 41 AND Y = 45 else
"100010011101" when X = 42 AND Y = 45 else
"100010011101" when X = 43 AND Y = 45 else
"100010011101" when X = 44 AND Y = 45 else
"100010011101" when X = 45 AND Y = 45 else
"100010011101" when X = 46 AND Y = 45 else
"100010011101" when X = 47 AND Y = 45 else
"100010011101" when X = 48 AND Y = 45 else
"100010011101" when X = 49 AND Y = 45 else
"110111011111" when X = 50 AND Y = 45 else
"110111011111" when X = 51 AND Y = 45 else
"110111011111" when X = 52 AND Y = 45 else
"110111011111" when X = 53 AND Y = 45 else
"110111011111" when X = 54 AND Y = 45 else
"110111011111" when X = 55 AND Y = 45 else
"110111011111" when X = 56 AND Y = 45 else
"110111011111" when X = 57 AND Y = 45 else
"110111011111" when X = 58 AND Y = 45 else
"110111011111" when X = 59 AND Y = 45 else
"111111111111" when X = 60 AND Y = 45 else
"111111111111" when X = 61 AND Y = 45 else
"111111111111" when X = 62 AND Y = 45 else
"111111111111" when X = 63 AND Y = 45 else
"111111111111" when X = 64 AND Y = 45 else
"111111111111" when X = 65 AND Y = 45 else
"111111111111" when X = 66 AND Y = 45 else
"111111111111" when X = 67 AND Y = 45 else
"111111111111" when X = 68 AND Y = 45 else
"111111111111" when X = 69 AND Y = 45 else
"111111111111" when X = 70 AND Y = 45 else
"111111111111" when X = 71 AND Y = 45 else
"111111111111" when X = 72 AND Y = 45 else
"111111111111" when X = 73 AND Y = 45 else
"111111111111" when X = 74 AND Y = 45 else
"111111111111" when X = 75 AND Y = 45 else
"111111111111" when X = 76 AND Y = 45 else
"111111111111" when X = 77 AND Y = 45 else
"111111111111" when X = 78 AND Y = 45 else
"111111111111" when X = 79 AND Y = 45 else
"111111111111" when X = 80 AND Y = 45 else
"111111111111" when X = 81 AND Y = 45 else
"111111111111" when X = 82 AND Y = 45 else
"111111111111" when X = 83 AND Y = 45 else
"111111111111" when X = 84 AND Y = 45 else
"111111111111" when X = 85 AND Y = 45 else
"111111111111" when X = 86 AND Y = 45 else
"111111111111" when X = 87 AND Y = 45 else
"111111111111" when X = 88 AND Y = 45 else
"111111111111" when X = 89 AND Y = 45 else
"111111111111" when X = 90 AND Y = 45 else
"111111111111" when X = 91 AND Y = 45 else
"111111111111" when X = 92 AND Y = 45 else
"111111111111" when X = 93 AND Y = 45 else
"111111111111" when X = 94 AND Y = 45 else
"111111111111" when X = 95 AND Y = 45 else
"111111111111" when X = 96 AND Y = 45 else
"111111111111" when X = 97 AND Y = 45 else
"111111111111" when X = 98 AND Y = 45 else
"111111111111" when X = 99 AND Y = 45 else
"111111111111" when X = 100 AND Y = 45 else
"111111111111" when X = 101 AND Y = 45 else
"111111111111" when X = 102 AND Y = 45 else
"111111111111" when X = 103 AND Y = 45 else
"111111111111" when X = 104 AND Y = 45 else
"111111111111" when X = 105 AND Y = 45 else
"111111111111" when X = 106 AND Y = 45 else
"111111111111" when X = 107 AND Y = 45 else
"111111111111" when X = 108 AND Y = 45 else
"111111111111" when X = 109 AND Y = 45 else
"111111111111" when X = 110 AND Y = 45 else
"111111111111" when X = 111 AND Y = 45 else
"111111111111" when X = 112 AND Y = 45 else
"111111111111" when X = 113 AND Y = 45 else
"111111111111" when X = 114 AND Y = 45 else
"111111111111" when X = 115 AND Y = 45 else
"111111111111" when X = 116 AND Y = 45 else
"111111111111" when X = 117 AND Y = 45 else
"111111111111" when X = 118 AND Y = 45 else
"111111111111" when X = 119 AND Y = 45 else
"111111111111" when X = 120 AND Y = 45 else
"111111111111" when X = 121 AND Y = 45 else
"111111111111" when X = 122 AND Y = 45 else
"111111111111" when X = 123 AND Y = 45 else
"111111111111" when X = 124 AND Y = 45 else
"111111111111" when X = 125 AND Y = 45 else
"111111111111" when X = 126 AND Y = 45 else
"111111111111" when X = 127 AND Y = 45 else
"111111111111" when X = 128 AND Y = 45 else
"111111111111" when X = 129 AND Y = 45 else
"111111111111" when X = 130 AND Y = 45 else
"111111111111" when X = 131 AND Y = 45 else
"111111111111" when X = 132 AND Y = 45 else
"111111111111" when X = 133 AND Y = 45 else
"111111111111" when X = 134 AND Y = 45 else
"111111111111" when X = 135 AND Y = 45 else
"111111111111" when X = 136 AND Y = 45 else
"111111111111" when X = 137 AND Y = 45 else
"111111111111" when X = 138 AND Y = 45 else
"111111111111" when X = 139 AND Y = 45 else
"111111111111" when X = 140 AND Y = 45 else
"111111111111" when X = 141 AND Y = 45 else
"111111111111" when X = 142 AND Y = 45 else
"111111111111" when X = 143 AND Y = 45 else
"111111111111" when X = 144 AND Y = 45 else
"111111111111" when X = 145 AND Y = 45 else
"111111111111" when X = 146 AND Y = 45 else
"111111111111" when X = 147 AND Y = 45 else
"111111111111" when X = 148 AND Y = 45 else
"111111111111" when X = 149 AND Y = 45 else
"111111111111" when X = 150 AND Y = 45 else
"111111111111" when X = 151 AND Y = 45 else
"111111111111" when X = 152 AND Y = 45 else
"111111111111" when X = 153 AND Y = 45 else
"111111111111" when X = 154 AND Y = 45 else
"111111111111" when X = 155 AND Y = 45 else
"111111111111" when X = 156 AND Y = 45 else
"111111111111" when X = 157 AND Y = 45 else
"111111111111" when X = 158 AND Y = 45 else
"111111111111" when X = 159 AND Y = 45 else
"111111111111" when X = 160 AND Y = 45 else
"111111111111" when X = 161 AND Y = 45 else
"111111111111" when X = 162 AND Y = 45 else
"111111111111" when X = 163 AND Y = 45 else
"111111111111" when X = 164 AND Y = 45 else
"111111111111" when X = 165 AND Y = 45 else
"111111111111" when X = 166 AND Y = 45 else
"111111111111" when X = 167 AND Y = 45 else
"111111111111" when X = 168 AND Y = 45 else
"111111111111" when X = 169 AND Y = 45 else
"111111111111" when X = 170 AND Y = 45 else
"111111111111" when X = 171 AND Y = 45 else
"111111111111" when X = 172 AND Y = 45 else
"111111111111" when X = 173 AND Y = 45 else
"111111111111" when X = 174 AND Y = 45 else
"111111111111" when X = 175 AND Y = 45 else
"111111111111" when X = 176 AND Y = 45 else
"111111111111" when X = 177 AND Y = 45 else
"111111111111" when X = 178 AND Y = 45 else
"111111111111" when X = 179 AND Y = 45 else
"111111111111" when X = 180 AND Y = 45 else
"111111111111" when X = 181 AND Y = 45 else
"111111111111" when X = 182 AND Y = 45 else
"111111111111" when X = 183 AND Y = 45 else
"111111111111" when X = 184 AND Y = 45 else
"111111111111" when X = 185 AND Y = 45 else
"111111111111" when X = 186 AND Y = 45 else
"111111111111" when X = 187 AND Y = 45 else
"111111111111" when X = 188 AND Y = 45 else
"111111111111" when X = 189 AND Y = 45 else
"111111111111" when X = 190 AND Y = 45 else
"111111111111" when X = 191 AND Y = 45 else
"111111111111" when X = 192 AND Y = 45 else
"111111111111" when X = 193 AND Y = 45 else
"111111111111" when X = 194 AND Y = 45 else
"111111111111" when X = 195 AND Y = 45 else
"111111111111" when X = 196 AND Y = 45 else
"111111111111" when X = 197 AND Y = 45 else
"111111111111" when X = 198 AND Y = 45 else
"111111111111" when X = 199 AND Y = 45 else
"111111111111" when X = 200 AND Y = 45 else
"111111111111" when X = 201 AND Y = 45 else
"111111111111" when X = 202 AND Y = 45 else
"111111111111" when X = 203 AND Y = 45 else
"111111111111" when X = 204 AND Y = 45 else
"111111111111" when X = 205 AND Y = 45 else
"111111111111" when X = 206 AND Y = 45 else
"111111111111" when X = 207 AND Y = 45 else
"111111111111" when X = 208 AND Y = 45 else
"111111111111" when X = 209 AND Y = 45 else
"111111111111" when X = 210 AND Y = 45 else
"111111111111" when X = 211 AND Y = 45 else
"111111111111" when X = 212 AND Y = 45 else
"111111111111" when X = 213 AND Y = 45 else
"111111111111" when X = 214 AND Y = 45 else
"111111111111" when X = 215 AND Y = 45 else
"111111111111" when X = 216 AND Y = 45 else
"111111111111" when X = 217 AND Y = 45 else
"111111111111" when X = 218 AND Y = 45 else
"111111111111" when X = 219 AND Y = 45 else
"111111111111" when X = 220 AND Y = 45 else
"111111111111" when X = 221 AND Y = 45 else
"111111111111" when X = 222 AND Y = 45 else
"111111111111" when X = 223 AND Y = 45 else
"111111111111" when X = 224 AND Y = 45 else
"111111111111" when X = 225 AND Y = 45 else
"111111111111" when X = 226 AND Y = 45 else
"111111111111" when X = 227 AND Y = 45 else
"111111111111" when X = 228 AND Y = 45 else
"111111111111" when X = 229 AND Y = 45 else
"111111111111" when X = 230 AND Y = 45 else
"111111111111" when X = 231 AND Y = 45 else
"111111111111" when X = 232 AND Y = 45 else
"111111111111" when X = 233 AND Y = 45 else
"111111111111" when X = 234 AND Y = 45 else
"111111111111" when X = 235 AND Y = 45 else
"111111111111" when X = 236 AND Y = 45 else
"111111111111" when X = 237 AND Y = 45 else
"111111111111" when X = 238 AND Y = 45 else
"111111111111" when X = 239 AND Y = 45 else
"111111111111" when X = 240 AND Y = 45 else
"111111111111" when X = 241 AND Y = 45 else
"111111111111" when X = 242 AND Y = 45 else
"111111111111" when X = 243 AND Y = 45 else
"111111111111" when X = 244 AND Y = 45 else
"111111111111" when X = 245 AND Y = 45 else
"111111111111" when X = 246 AND Y = 45 else
"111111111111" when X = 247 AND Y = 45 else
"111111111111" when X = 248 AND Y = 45 else
"111111111111" when X = 249 AND Y = 45 else
"111111111111" when X = 250 AND Y = 45 else
"111111111111" when X = 251 AND Y = 45 else
"111111111111" when X = 252 AND Y = 45 else
"111111111111" when X = 253 AND Y = 45 else
"111111111111" when X = 254 AND Y = 45 else
"111111111111" when X = 255 AND Y = 45 else
"111111111111" when X = 256 AND Y = 45 else
"111111111111" when X = 257 AND Y = 45 else
"111111111111" when X = 258 AND Y = 45 else
"111111111111" when X = 259 AND Y = 45 else
"111111111111" when X = 260 AND Y = 45 else
"111111111111" when X = 261 AND Y = 45 else
"111111111111" when X = 262 AND Y = 45 else
"111111111111" when X = 263 AND Y = 45 else
"111111111111" when X = 264 AND Y = 45 else
"110111011111" when X = 265 AND Y = 45 else
"110111011111" when X = 266 AND Y = 45 else
"110111011111" when X = 267 AND Y = 45 else
"110111011111" when X = 268 AND Y = 45 else
"110111011111" when X = 269 AND Y = 45 else
"110111011111" when X = 270 AND Y = 45 else
"110111011111" when X = 271 AND Y = 45 else
"110111011111" when X = 272 AND Y = 45 else
"110111011111" when X = 273 AND Y = 45 else
"110111011111" when X = 274 AND Y = 45 else
"110111011111" when X = 275 AND Y = 45 else
"110111011111" when X = 276 AND Y = 45 else
"110111011111" when X = 277 AND Y = 45 else
"110111011111" when X = 278 AND Y = 45 else
"110111011111" when X = 279 AND Y = 45 else
"000000000000" when X = 280 AND Y = 45 else
"000000000000" when X = 281 AND Y = 45 else
"000000000000" when X = 282 AND Y = 45 else
"000000000000" when X = 283 AND Y = 45 else
"000000000000" when X = 284 AND Y = 45 else
"000000000000" when X = 285 AND Y = 45 else
"000000000000" when X = 286 AND Y = 45 else
"000000000000" when X = 287 AND Y = 45 else
"000000000000" when X = 288 AND Y = 45 else
"000000000000" when X = 289 AND Y = 45 else
"000000000000" when X = 290 AND Y = 45 else
"000000000000" when X = 291 AND Y = 45 else
"000000000000" when X = 292 AND Y = 45 else
"000000000000" when X = 293 AND Y = 45 else
"000000000000" when X = 294 AND Y = 45 else
"000000000000" when X = 295 AND Y = 45 else
"000000000000" when X = 296 AND Y = 45 else
"000000000000" when X = 297 AND Y = 45 else
"000000000000" when X = 298 AND Y = 45 else
"000000000000" when X = 299 AND Y = 45 else
"000000000000" when X = 300 AND Y = 45 else
"000000000000" when X = 301 AND Y = 45 else
"000000000000" when X = 302 AND Y = 45 else
"000000000000" when X = 303 AND Y = 45 else
"000000000000" when X = 304 AND Y = 45 else
"000000000000" when X = 305 AND Y = 45 else
"000000000000" when X = 306 AND Y = 45 else
"000000000000" when X = 307 AND Y = 45 else
"000000000000" when X = 308 AND Y = 45 else
"000000000000" when X = 309 AND Y = 45 else
"000000000000" when X = 310 AND Y = 45 else
"000000000000" when X = 311 AND Y = 45 else
"000000000000" when X = 312 AND Y = 45 else
"000000000000" when X = 313 AND Y = 45 else
"000000000000" when X = 314 AND Y = 45 else
"000000000000" when X = 315 AND Y = 45 else
"000000000000" when X = 316 AND Y = 45 else
"000000000000" when X = 317 AND Y = 45 else
"000000000000" when X = 318 AND Y = 45 else
"000000000000" when X = 319 AND Y = 45 else
"000000000000" when X = 320 AND Y = 45 else
"000000000000" when X = 321 AND Y = 45 else
"000000000000" when X = 322 AND Y = 45 else
"000000000000" when X = 323 AND Y = 45 else
"000000000000" when X = 324 AND Y = 45 else
"000000000000" when X = 0 AND Y = 46 else
"000000000000" when X = 1 AND Y = 46 else
"000000000000" when X = 2 AND Y = 46 else
"000000000000" when X = 3 AND Y = 46 else
"000000000000" when X = 4 AND Y = 46 else
"000000000000" when X = 5 AND Y = 46 else
"000000000000" when X = 6 AND Y = 46 else
"000000000000" when X = 7 AND Y = 46 else
"000000000000" when X = 8 AND Y = 46 else
"000000000000" when X = 9 AND Y = 46 else
"000000000000" when X = 10 AND Y = 46 else
"000000000000" when X = 11 AND Y = 46 else
"000000000000" when X = 12 AND Y = 46 else
"000000000000" when X = 13 AND Y = 46 else
"000000000000" when X = 14 AND Y = 46 else
"000000000000" when X = 15 AND Y = 46 else
"000000000000" when X = 16 AND Y = 46 else
"000000000000" when X = 17 AND Y = 46 else
"000000000000" when X = 18 AND Y = 46 else
"000000000000" when X = 19 AND Y = 46 else
"000000000000" when X = 20 AND Y = 46 else
"000000000000" when X = 21 AND Y = 46 else
"000000000000" when X = 22 AND Y = 46 else
"000000000000" when X = 23 AND Y = 46 else
"000000000000" when X = 24 AND Y = 46 else
"000000000000" when X = 25 AND Y = 46 else
"000000000000" when X = 26 AND Y = 46 else
"000000000000" when X = 27 AND Y = 46 else
"000000000000" when X = 28 AND Y = 46 else
"000000000000" when X = 29 AND Y = 46 else
"000000000000" when X = 30 AND Y = 46 else
"000000000000" when X = 31 AND Y = 46 else
"000000000000" when X = 32 AND Y = 46 else
"000000000000" when X = 33 AND Y = 46 else
"000000000000" when X = 34 AND Y = 46 else
"000000000000" when X = 35 AND Y = 46 else
"000000000000" when X = 36 AND Y = 46 else
"000000000000" when X = 37 AND Y = 46 else
"000000000000" when X = 38 AND Y = 46 else
"000000000000" when X = 39 AND Y = 46 else
"100010011101" when X = 40 AND Y = 46 else
"100010011101" when X = 41 AND Y = 46 else
"100010011101" when X = 42 AND Y = 46 else
"100010011101" when X = 43 AND Y = 46 else
"100010011101" when X = 44 AND Y = 46 else
"100010011101" when X = 45 AND Y = 46 else
"100010011101" when X = 46 AND Y = 46 else
"100010011101" when X = 47 AND Y = 46 else
"100010011101" when X = 48 AND Y = 46 else
"100010011101" when X = 49 AND Y = 46 else
"110111011111" when X = 50 AND Y = 46 else
"110111011111" when X = 51 AND Y = 46 else
"110111011111" when X = 52 AND Y = 46 else
"110111011111" when X = 53 AND Y = 46 else
"110111011111" when X = 54 AND Y = 46 else
"110111011111" when X = 55 AND Y = 46 else
"110111011111" when X = 56 AND Y = 46 else
"110111011111" when X = 57 AND Y = 46 else
"110111011111" when X = 58 AND Y = 46 else
"110111011111" when X = 59 AND Y = 46 else
"111111111111" when X = 60 AND Y = 46 else
"111111111111" when X = 61 AND Y = 46 else
"111111111111" when X = 62 AND Y = 46 else
"111111111111" when X = 63 AND Y = 46 else
"111111111111" when X = 64 AND Y = 46 else
"111111111111" when X = 65 AND Y = 46 else
"111111111111" when X = 66 AND Y = 46 else
"111111111111" when X = 67 AND Y = 46 else
"111111111111" when X = 68 AND Y = 46 else
"111111111111" when X = 69 AND Y = 46 else
"111111111111" when X = 70 AND Y = 46 else
"111111111111" when X = 71 AND Y = 46 else
"111111111111" when X = 72 AND Y = 46 else
"111111111111" when X = 73 AND Y = 46 else
"111111111111" when X = 74 AND Y = 46 else
"111111111111" when X = 75 AND Y = 46 else
"111111111111" when X = 76 AND Y = 46 else
"111111111111" when X = 77 AND Y = 46 else
"111111111111" when X = 78 AND Y = 46 else
"111111111111" when X = 79 AND Y = 46 else
"111111111111" when X = 80 AND Y = 46 else
"111111111111" when X = 81 AND Y = 46 else
"111111111111" when X = 82 AND Y = 46 else
"111111111111" when X = 83 AND Y = 46 else
"111111111111" when X = 84 AND Y = 46 else
"111111111111" when X = 85 AND Y = 46 else
"111111111111" when X = 86 AND Y = 46 else
"111111111111" when X = 87 AND Y = 46 else
"111111111111" when X = 88 AND Y = 46 else
"111111111111" when X = 89 AND Y = 46 else
"111111111111" when X = 90 AND Y = 46 else
"111111111111" when X = 91 AND Y = 46 else
"111111111111" when X = 92 AND Y = 46 else
"111111111111" when X = 93 AND Y = 46 else
"111111111111" when X = 94 AND Y = 46 else
"111111111111" when X = 95 AND Y = 46 else
"111111111111" when X = 96 AND Y = 46 else
"111111111111" when X = 97 AND Y = 46 else
"111111111111" when X = 98 AND Y = 46 else
"111111111111" when X = 99 AND Y = 46 else
"111111111111" when X = 100 AND Y = 46 else
"111111111111" when X = 101 AND Y = 46 else
"111111111111" when X = 102 AND Y = 46 else
"111111111111" when X = 103 AND Y = 46 else
"111111111111" when X = 104 AND Y = 46 else
"111111111111" when X = 105 AND Y = 46 else
"111111111111" when X = 106 AND Y = 46 else
"111111111111" when X = 107 AND Y = 46 else
"111111111111" when X = 108 AND Y = 46 else
"111111111111" when X = 109 AND Y = 46 else
"111111111111" when X = 110 AND Y = 46 else
"111111111111" when X = 111 AND Y = 46 else
"111111111111" when X = 112 AND Y = 46 else
"111111111111" when X = 113 AND Y = 46 else
"111111111111" when X = 114 AND Y = 46 else
"111111111111" when X = 115 AND Y = 46 else
"111111111111" when X = 116 AND Y = 46 else
"111111111111" when X = 117 AND Y = 46 else
"111111111111" when X = 118 AND Y = 46 else
"111111111111" when X = 119 AND Y = 46 else
"111111111111" when X = 120 AND Y = 46 else
"111111111111" when X = 121 AND Y = 46 else
"111111111111" when X = 122 AND Y = 46 else
"111111111111" when X = 123 AND Y = 46 else
"111111111111" when X = 124 AND Y = 46 else
"111111111111" when X = 125 AND Y = 46 else
"111111111111" when X = 126 AND Y = 46 else
"111111111111" when X = 127 AND Y = 46 else
"111111111111" when X = 128 AND Y = 46 else
"111111111111" when X = 129 AND Y = 46 else
"111111111111" when X = 130 AND Y = 46 else
"111111111111" when X = 131 AND Y = 46 else
"111111111111" when X = 132 AND Y = 46 else
"111111111111" when X = 133 AND Y = 46 else
"111111111111" when X = 134 AND Y = 46 else
"111111111111" when X = 135 AND Y = 46 else
"111111111111" when X = 136 AND Y = 46 else
"111111111111" when X = 137 AND Y = 46 else
"111111111111" when X = 138 AND Y = 46 else
"111111111111" when X = 139 AND Y = 46 else
"111111111111" when X = 140 AND Y = 46 else
"111111111111" when X = 141 AND Y = 46 else
"111111111111" when X = 142 AND Y = 46 else
"111111111111" when X = 143 AND Y = 46 else
"111111111111" when X = 144 AND Y = 46 else
"111111111111" when X = 145 AND Y = 46 else
"111111111111" when X = 146 AND Y = 46 else
"111111111111" when X = 147 AND Y = 46 else
"111111111111" when X = 148 AND Y = 46 else
"111111111111" when X = 149 AND Y = 46 else
"111111111111" when X = 150 AND Y = 46 else
"111111111111" when X = 151 AND Y = 46 else
"111111111111" when X = 152 AND Y = 46 else
"111111111111" when X = 153 AND Y = 46 else
"111111111111" when X = 154 AND Y = 46 else
"111111111111" when X = 155 AND Y = 46 else
"111111111111" when X = 156 AND Y = 46 else
"111111111111" when X = 157 AND Y = 46 else
"111111111111" when X = 158 AND Y = 46 else
"111111111111" when X = 159 AND Y = 46 else
"111111111111" when X = 160 AND Y = 46 else
"111111111111" when X = 161 AND Y = 46 else
"111111111111" when X = 162 AND Y = 46 else
"111111111111" when X = 163 AND Y = 46 else
"111111111111" when X = 164 AND Y = 46 else
"111111111111" when X = 165 AND Y = 46 else
"111111111111" when X = 166 AND Y = 46 else
"111111111111" when X = 167 AND Y = 46 else
"111111111111" when X = 168 AND Y = 46 else
"111111111111" when X = 169 AND Y = 46 else
"111111111111" when X = 170 AND Y = 46 else
"111111111111" when X = 171 AND Y = 46 else
"111111111111" when X = 172 AND Y = 46 else
"111111111111" when X = 173 AND Y = 46 else
"111111111111" when X = 174 AND Y = 46 else
"111111111111" when X = 175 AND Y = 46 else
"111111111111" when X = 176 AND Y = 46 else
"111111111111" when X = 177 AND Y = 46 else
"111111111111" when X = 178 AND Y = 46 else
"111111111111" when X = 179 AND Y = 46 else
"111111111111" when X = 180 AND Y = 46 else
"111111111111" when X = 181 AND Y = 46 else
"111111111111" when X = 182 AND Y = 46 else
"111111111111" when X = 183 AND Y = 46 else
"111111111111" when X = 184 AND Y = 46 else
"111111111111" when X = 185 AND Y = 46 else
"111111111111" when X = 186 AND Y = 46 else
"111111111111" when X = 187 AND Y = 46 else
"111111111111" when X = 188 AND Y = 46 else
"111111111111" when X = 189 AND Y = 46 else
"111111111111" when X = 190 AND Y = 46 else
"111111111111" when X = 191 AND Y = 46 else
"111111111111" when X = 192 AND Y = 46 else
"111111111111" when X = 193 AND Y = 46 else
"111111111111" when X = 194 AND Y = 46 else
"111111111111" when X = 195 AND Y = 46 else
"111111111111" when X = 196 AND Y = 46 else
"111111111111" when X = 197 AND Y = 46 else
"111111111111" when X = 198 AND Y = 46 else
"111111111111" when X = 199 AND Y = 46 else
"111111111111" when X = 200 AND Y = 46 else
"111111111111" when X = 201 AND Y = 46 else
"111111111111" when X = 202 AND Y = 46 else
"111111111111" when X = 203 AND Y = 46 else
"111111111111" when X = 204 AND Y = 46 else
"111111111111" when X = 205 AND Y = 46 else
"111111111111" when X = 206 AND Y = 46 else
"111111111111" when X = 207 AND Y = 46 else
"111111111111" when X = 208 AND Y = 46 else
"111111111111" when X = 209 AND Y = 46 else
"111111111111" when X = 210 AND Y = 46 else
"111111111111" when X = 211 AND Y = 46 else
"111111111111" when X = 212 AND Y = 46 else
"111111111111" when X = 213 AND Y = 46 else
"111111111111" when X = 214 AND Y = 46 else
"111111111111" when X = 215 AND Y = 46 else
"111111111111" when X = 216 AND Y = 46 else
"111111111111" when X = 217 AND Y = 46 else
"111111111111" when X = 218 AND Y = 46 else
"111111111111" when X = 219 AND Y = 46 else
"111111111111" when X = 220 AND Y = 46 else
"111111111111" when X = 221 AND Y = 46 else
"111111111111" when X = 222 AND Y = 46 else
"111111111111" when X = 223 AND Y = 46 else
"111111111111" when X = 224 AND Y = 46 else
"111111111111" when X = 225 AND Y = 46 else
"111111111111" when X = 226 AND Y = 46 else
"111111111111" when X = 227 AND Y = 46 else
"111111111111" when X = 228 AND Y = 46 else
"111111111111" when X = 229 AND Y = 46 else
"111111111111" when X = 230 AND Y = 46 else
"111111111111" when X = 231 AND Y = 46 else
"111111111111" when X = 232 AND Y = 46 else
"111111111111" when X = 233 AND Y = 46 else
"111111111111" when X = 234 AND Y = 46 else
"111111111111" when X = 235 AND Y = 46 else
"111111111111" when X = 236 AND Y = 46 else
"111111111111" when X = 237 AND Y = 46 else
"111111111111" when X = 238 AND Y = 46 else
"111111111111" when X = 239 AND Y = 46 else
"111111111111" when X = 240 AND Y = 46 else
"111111111111" when X = 241 AND Y = 46 else
"111111111111" when X = 242 AND Y = 46 else
"111111111111" when X = 243 AND Y = 46 else
"111111111111" when X = 244 AND Y = 46 else
"111111111111" when X = 245 AND Y = 46 else
"111111111111" when X = 246 AND Y = 46 else
"111111111111" when X = 247 AND Y = 46 else
"111111111111" when X = 248 AND Y = 46 else
"111111111111" when X = 249 AND Y = 46 else
"111111111111" when X = 250 AND Y = 46 else
"111111111111" when X = 251 AND Y = 46 else
"111111111111" when X = 252 AND Y = 46 else
"111111111111" when X = 253 AND Y = 46 else
"111111111111" when X = 254 AND Y = 46 else
"111111111111" when X = 255 AND Y = 46 else
"111111111111" when X = 256 AND Y = 46 else
"111111111111" when X = 257 AND Y = 46 else
"111111111111" when X = 258 AND Y = 46 else
"111111111111" when X = 259 AND Y = 46 else
"111111111111" when X = 260 AND Y = 46 else
"111111111111" when X = 261 AND Y = 46 else
"111111111111" when X = 262 AND Y = 46 else
"111111111111" when X = 263 AND Y = 46 else
"111111111111" when X = 264 AND Y = 46 else
"110111011111" when X = 265 AND Y = 46 else
"110111011111" when X = 266 AND Y = 46 else
"110111011111" when X = 267 AND Y = 46 else
"110111011111" when X = 268 AND Y = 46 else
"110111011111" when X = 269 AND Y = 46 else
"110111011111" when X = 270 AND Y = 46 else
"110111011111" when X = 271 AND Y = 46 else
"110111011111" when X = 272 AND Y = 46 else
"110111011111" when X = 273 AND Y = 46 else
"110111011111" when X = 274 AND Y = 46 else
"110111011111" when X = 275 AND Y = 46 else
"110111011111" when X = 276 AND Y = 46 else
"110111011111" when X = 277 AND Y = 46 else
"110111011111" when X = 278 AND Y = 46 else
"110111011111" when X = 279 AND Y = 46 else
"000000000000" when X = 280 AND Y = 46 else
"000000000000" when X = 281 AND Y = 46 else
"000000000000" when X = 282 AND Y = 46 else
"000000000000" when X = 283 AND Y = 46 else
"000000000000" when X = 284 AND Y = 46 else
"000000000000" when X = 285 AND Y = 46 else
"000000000000" when X = 286 AND Y = 46 else
"000000000000" when X = 287 AND Y = 46 else
"000000000000" when X = 288 AND Y = 46 else
"000000000000" when X = 289 AND Y = 46 else
"000000000000" when X = 290 AND Y = 46 else
"000000000000" when X = 291 AND Y = 46 else
"000000000000" when X = 292 AND Y = 46 else
"000000000000" when X = 293 AND Y = 46 else
"000000000000" when X = 294 AND Y = 46 else
"000000000000" when X = 295 AND Y = 46 else
"000000000000" when X = 296 AND Y = 46 else
"000000000000" when X = 297 AND Y = 46 else
"000000000000" when X = 298 AND Y = 46 else
"000000000000" when X = 299 AND Y = 46 else
"000000000000" when X = 300 AND Y = 46 else
"000000000000" when X = 301 AND Y = 46 else
"000000000000" when X = 302 AND Y = 46 else
"000000000000" when X = 303 AND Y = 46 else
"000000000000" when X = 304 AND Y = 46 else
"000000000000" when X = 305 AND Y = 46 else
"000000000000" when X = 306 AND Y = 46 else
"000000000000" when X = 307 AND Y = 46 else
"000000000000" when X = 308 AND Y = 46 else
"000000000000" when X = 309 AND Y = 46 else
"000000000000" when X = 310 AND Y = 46 else
"000000000000" when X = 311 AND Y = 46 else
"000000000000" when X = 312 AND Y = 46 else
"000000000000" when X = 313 AND Y = 46 else
"000000000000" when X = 314 AND Y = 46 else
"000000000000" when X = 315 AND Y = 46 else
"000000000000" when X = 316 AND Y = 46 else
"000000000000" when X = 317 AND Y = 46 else
"000000000000" when X = 318 AND Y = 46 else
"000000000000" when X = 319 AND Y = 46 else
"000000000000" when X = 320 AND Y = 46 else
"000000000000" when X = 321 AND Y = 46 else
"000000000000" when X = 322 AND Y = 46 else
"000000000000" when X = 323 AND Y = 46 else
"000000000000" when X = 324 AND Y = 46 else
"000000000000" when X = 0 AND Y = 47 else
"000000000000" when X = 1 AND Y = 47 else
"000000000000" when X = 2 AND Y = 47 else
"000000000000" when X = 3 AND Y = 47 else
"000000000000" when X = 4 AND Y = 47 else
"000000000000" when X = 5 AND Y = 47 else
"000000000000" when X = 6 AND Y = 47 else
"000000000000" when X = 7 AND Y = 47 else
"000000000000" when X = 8 AND Y = 47 else
"000000000000" when X = 9 AND Y = 47 else
"000000000000" when X = 10 AND Y = 47 else
"000000000000" when X = 11 AND Y = 47 else
"000000000000" when X = 12 AND Y = 47 else
"000000000000" when X = 13 AND Y = 47 else
"000000000000" when X = 14 AND Y = 47 else
"000000000000" when X = 15 AND Y = 47 else
"000000000000" when X = 16 AND Y = 47 else
"000000000000" when X = 17 AND Y = 47 else
"000000000000" when X = 18 AND Y = 47 else
"000000000000" when X = 19 AND Y = 47 else
"000000000000" when X = 20 AND Y = 47 else
"000000000000" when X = 21 AND Y = 47 else
"000000000000" when X = 22 AND Y = 47 else
"000000000000" when X = 23 AND Y = 47 else
"000000000000" when X = 24 AND Y = 47 else
"000000000000" when X = 25 AND Y = 47 else
"000000000000" when X = 26 AND Y = 47 else
"000000000000" when X = 27 AND Y = 47 else
"000000000000" when X = 28 AND Y = 47 else
"000000000000" when X = 29 AND Y = 47 else
"000000000000" when X = 30 AND Y = 47 else
"000000000000" when X = 31 AND Y = 47 else
"000000000000" when X = 32 AND Y = 47 else
"000000000000" when X = 33 AND Y = 47 else
"000000000000" when X = 34 AND Y = 47 else
"000000000000" when X = 35 AND Y = 47 else
"000000000000" when X = 36 AND Y = 47 else
"000000000000" when X = 37 AND Y = 47 else
"000000000000" when X = 38 AND Y = 47 else
"000000000000" when X = 39 AND Y = 47 else
"100010011101" when X = 40 AND Y = 47 else
"100010011101" when X = 41 AND Y = 47 else
"100010011101" when X = 42 AND Y = 47 else
"100010011101" when X = 43 AND Y = 47 else
"100010011101" when X = 44 AND Y = 47 else
"100010011101" when X = 45 AND Y = 47 else
"100010011101" when X = 46 AND Y = 47 else
"100010011101" when X = 47 AND Y = 47 else
"100010011101" when X = 48 AND Y = 47 else
"100010011101" when X = 49 AND Y = 47 else
"110111011111" when X = 50 AND Y = 47 else
"110111011111" when X = 51 AND Y = 47 else
"110111011111" when X = 52 AND Y = 47 else
"110111011111" when X = 53 AND Y = 47 else
"110111011111" when X = 54 AND Y = 47 else
"110111011111" when X = 55 AND Y = 47 else
"110111011111" when X = 56 AND Y = 47 else
"110111011111" when X = 57 AND Y = 47 else
"110111011111" when X = 58 AND Y = 47 else
"110111011111" when X = 59 AND Y = 47 else
"111111111111" when X = 60 AND Y = 47 else
"111111111111" when X = 61 AND Y = 47 else
"111111111111" when X = 62 AND Y = 47 else
"111111111111" when X = 63 AND Y = 47 else
"111111111111" when X = 64 AND Y = 47 else
"111111111111" when X = 65 AND Y = 47 else
"111111111111" when X = 66 AND Y = 47 else
"111111111111" when X = 67 AND Y = 47 else
"111111111111" when X = 68 AND Y = 47 else
"111111111111" when X = 69 AND Y = 47 else
"111111111111" when X = 70 AND Y = 47 else
"111111111111" when X = 71 AND Y = 47 else
"111111111111" when X = 72 AND Y = 47 else
"111111111111" when X = 73 AND Y = 47 else
"111111111111" when X = 74 AND Y = 47 else
"111111111111" when X = 75 AND Y = 47 else
"111111111111" when X = 76 AND Y = 47 else
"111111111111" when X = 77 AND Y = 47 else
"111111111111" when X = 78 AND Y = 47 else
"111111111111" when X = 79 AND Y = 47 else
"111111111111" when X = 80 AND Y = 47 else
"111111111111" when X = 81 AND Y = 47 else
"111111111111" when X = 82 AND Y = 47 else
"111111111111" when X = 83 AND Y = 47 else
"111111111111" when X = 84 AND Y = 47 else
"111111111111" when X = 85 AND Y = 47 else
"111111111111" when X = 86 AND Y = 47 else
"111111111111" when X = 87 AND Y = 47 else
"111111111111" when X = 88 AND Y = 47 else
"111111111111" when X = 89 AND Y = 47 else
"111111111111" when X = 90 AND Y = 47 else
"111111111111" when X = 91 AND Y = 47 else
"111111111111" when X = 92 AND Y = 47 else
"111111111111" when X = 93 AND Y = 47 else
"111111111111" when X = 94 AND Y = 47 else
"111111111111" when X = 95 AND Y = 47 else
"111111111111" when X = 96 AND Y = 47 else
"111111111111" when X = 97 AND Y = 47 else
"111111111111" when X = 98 AND Y = 47 else
"111111111111" when X = 99 AND Y = 47 else
"111111111111" when X = 100 AND Y = 47 else
"111111111111" when X = 101 AND Y = 47 else
"111111111111" when X = 102 AND Y = 47 else
"111111111111" when X = 103 AND Y = 47 else
"111111111111" when X = 104 AND Y = 47 else
"111111111111" when X = 105 AND Y = 47 else
"111111111111" when X = 106 AND Y = 47 else
"111111111111" when X = 107 AND Y = 47 else
"111111111111" when X = 108 AND Y = 47 else
"111111111111" when X = 109 AND Y = 47 else
"111111111111" when X = 110 AND Y = 47 else
"111111111111" when X = 111 AND Y = 47 else
"111111111111" when X = 112 AND Y = 47 else
"111111111111" when X = 113 AND Y = 47 else
"111111111111" when X = 114 AND Y = 47 else
"111111111111" when X = 115 AND Y = 47 else
"111111111111" when X = 116 AND Y = 47 else
"111111111111" when X = 117 AND Y = 47 else
"111111111111" when X = 118 AND Y = 47 else
"111111111111" when X = 119 AND Y = 47 else
"111111111111" when X = 120 AND Y = 47 else
"111111111111" when X = 121 AND Y = 47 else
"111111111111" when X = 122 AND Y = 47 else
"111111111111" when X = 123 AND Y = 47 else
"111111111111" when X = 124 AND Y = 47 else
"111111111111" when X = 125 AND Y = 47 else
"111111111111" when X = 126 AND Y = 47 else
"111111111111" when X = 127 AND Y = 47 else
"111111111111" when X = 128 AND Y = 47 else
"111111111111" when X = 129 AND Y = 47 else
"111111111111" when X = 130 AND Y = 47 else
"111111111111" when X = 131 AND Y = 47 else
"111111111111" when X = 132 AND Y = 47 else
"111111111111" when X = 133 AND Y = 47 else
"111111111111" when X = 134 AND Y = 47 else
"111111111111" when X = 135 AND Y = 47 else
"111111111111" when X = 136 AND Y = 47 else
"111111111111" when X = 137 AND Y = 47 else
"111111111111" when X = 138 AND Y = 47 else
"111111111111" when X = 139 AND Y = 47 else
"111111111111" when X = 140 AND Y = 47 else
"111111111111" when X = 141 AND Y = 47 else
"111111111111" when X = 142 AND Y = 47 else
"111111111111" when X = 143 AND Y = 47 else
"111111111111" when X = 144 AND Y = 47 else
"111111111111" when X = 145 AND Y = 47 else
"111111111111" when X = 146 AND Y = 47 else
"111111111111" when X = 147 AND Y = 47 else
"111111111111" when X = 148 AND Y = 47 else
"111111111111" when X = 149 AND Y = 47 else
"111111111111" when X = 150 AND Y = 47 else
"111111111111" when X = 151 AND Y = 47 else
"111111111111" when X = 152 AND Y = 47 else
"111111111111" when X = 153 AND Y = 47 else
"111111111111" when X = 154 AND Y = 47 else
"111111111111" when X = 155 AND Y = 47 else
"111111111111" when X = 156 AND Y = 47 else
"111111111111" when X = 157 AND Y = 47 else
"111111111111" when X = 158 AND Y = 47 else
"111111111111" when X = 159 AND Y = 47 else
"111111111111" when X = 160 AND Y = 47 else
"111111111111" when X = 161 AND Y = 47 else
"111111111111" when X = 162 AND Y = 47 else
"111111111111" when X = 163 AND Y = 47 else
"111111111111" when X = 164 AND Y = 47 else
"111111111111" when X = 165 AND Y = 47 else
"111111111111" when X = 166 AND Y = 47 else
"111111111111" when X = 167 AND Y = 47 else
"111111111111" when X = 168 AND Y = 47 else
"111111111111" when X = 169 AND Y = 47 else
"111111111111" when X = 170 AND Y = 47 else
"111111111111" when X = 171 AND Y = 47 else
"111111111111" when X = 172 AND Y = 47 else
"111111111111" when X = 173 AND Y = 47 else
"111111111111" when X = 174 AND Y = 47 else
"111111111111" when X = 175 AND Y = 47 else
"111111111111" when X = 176 AND Y = 47 else
"111111111111" when X = 177 AND Y = 47 else
"111111111111" when X = 178 AND Y = 47 else
"111111111111" when X = 179 AND Y = 47 else
"111111111111" when X = 180 AND Y = 47 else
"111111111111" when X = 181 AND Y = 47 else
"111111111111" when X = 182 AND Y = 47 else
"111111111111" when X = 183 AND Y = 47 else
"111111111111" when X = 184 AND Y = 47 else
"111111111111" when X = 185 AND Y = 47 else
"111111111111" when X = 186 AND Y = 47 else
"111111111111" when X = 187 AND Y = 47 else
"111111111111" when X = 188 AND Y = 47 else
"111111111111" when X = 189 AND Y = 47 else
"111111111111" when X = 190 AND Y = 47 else
"111111111111" when X = 191 AND Y = 47 else
"111111111111" when X = 192 AND Y = 47 else
"111111111111" when X = 193 AND Y = 47 else
"111111111111" when X = 194 AND Y = 47 else
"111111111111" when X = 195 AND Y = 47 else
"111111111111" when X = 196 AND Y = 47 else
"111111111111" when X = 197 AND Y = 47 else
"111111111111" when X = 198 AND Y = 47 else
"111111111111" when X = 199 AND Y = 47 else
"111111111111" when X = 200 AND Y = 47 else
"111111111111" when X = 201 AND Y = 47 else
"111111111111" when X = 202 AND Y = 47 else
"111111111111" when X = 203 AND Y = 47 else
"111111111111" when X = 204 AND Y = 47 else
"111111111111" when X = 205 AND Y = 47 else
"111111111111" when X = 206 AND Y = 47 else
"111111111111" when X = 207 AND Y = 47 else
"111111111111" when X = 208 AND Y = 47 else
"111111111111" when X = 209 AND Y = 47 else
"111111111111" when X = 210 AND Y = 47 else
"111111111111" when X = 211 AND Y = 47 else
"111111111111" when X = 212 AND Y = 47 else
"111111111111" when X = 213 AND Y = 47 else
"111111111111" when X = 214 AND Y = 47 else
"111111111111" when X = 215 AND Y = 47 else
"111111111111" when X = 216 AND Y = 47 else
"111111111111" when X = 217 AND Y = 47 else
"111111111111" when X = 218 AND Y = 47 else
"111111111111" when X = 219 AND Y = 47 else
"111111111111" when X = 220 AND Y = 47 else
"111111111111" when X = 221 AND Y = 47 else
"111111111111" when X = 222 AND Y = 47 else
"111111111111" when X = 223 AND Y = 47 else
"111111111111" when X = 224 AND Y = 47 else
"111111111111" when X = 225 AND Y = 47 else
"111111111111" when X = 226 AND Y = 47 else
"111111111111" when X = 227 AND Y = 47 else
"111111111111" when X = 228 AND Y = 47 else
"111111111111" when X = 229 AND Y = 47 else
"111111111111" when X = 230 AND Y = 47 else
"111111111111" when X = 231 AND Y = 47 else
"111111111111" when X = 232 AND Y = 47 else
"111111111111" when X = 233 AND Y = 47 else
"111111111111" when X = 234 AND Y = 47 else
"111111111111" when X = 235 AND Y = 47 else
"111111111111" when X = 236 AND Y = 47 else
"111111111111" when X = 237 AND Y = 47 else
"111111111111" when X = 238 AND Y = 47 else
"111111111111" when X = 239 AND Y = 47 else
"111111111111" when X = 240 AND Y = 47 else
"111111111111" when X = 241 AND Y = 47 else
"111111111111" when X = 242 AND Y = 47 else
"111111111111" when X = 243 AND Y = 47 else
"111111111111" when X = 244 AND Y = 47 else
"111111111111" when X = 245 AND Y = 47 else
"111111111111" when X = 246 AND Y = 47 else
"111111111111" when X = 247 AND Y = 47 else
"111111111111" when X = 248 AND Y = 47 else
"111111111111" when X = 249 AND Y = 47 else
"111111111111" when X = 250 AND Y = 47 else
"111111111111" when X = 251 AND Y = 47 else
"111111111111" when X = 252 AND Y = 47 else
"111111111111" when X = 253 AND Y = 47 else
"111111111111" when X = 254 AND Y = 47 else
"111111111111" when X = 255 AND Y = 47 else
"111111111111" when X = 256 AND Y = 47 else
"111111111111" when X = 257 AND Y = 47 else
"111111111111" when X = 258 AND Y = 47 else
"111111111111" when X = 259 AND Y = 47 else
"111111111111" when X = 260 AND Y = 47 else
"111111111111" when X = 261 AND Y = 47 else
"111111111111" when X = 262 AND Y = 47 else
"111111111111" when X = 263 AND Y = 47 else
"111111111111" when X = 264 AND Y = 47 else
"110111011111" when X = 265 AND Y = 47 else
"110111011111" when X = 266 AND Y = 47 else
"110111011111" when X = 267 AND Y = 47 else
"110111011111" when X = 268 AND Y = 47 else
"110111011111" when X = 269 AND Y = 47 else
"110111011111" when X = 270 AND Y = 47 else
"110111011111" when X = 271 AND Y = 47 else
"110111011111" when X = 272 AND Y = 47 else
"110111011111" when X = 273 AND Y = 47 else
"110111011111" when X = 274 AND Y = 47 else
"110111011111" when X = 275 AND Y = 47 else
"110111011111" when X = 276 AND Y = 47 else
"110111011111" when X = 277 AND Y = 47 else
"110111011111" when X = 278 AND Y = 47 else
"110111011111" when X = 279 AND Y = 47 else
"000000000000" when X = 280 AND Y = 47 else
"000000000000" when X = 281 AND Y = 47 else
"000000000000" when X = 282 AND Y = 47 else
"000000000000" when X = 283 AND Y = 47 else
"000000000000" when X = 284 AND Y = 47 else
"000000000000" when X = 285 AND Y = 47 else
"000000000000" when X = 286 AND Y = 47 else
"000000000000" when X = 287 AND Y = 47 else
"000000000000" when X = 288 AND Y = 47 else
"000000000000" when X = 289 AND Y = 47 else
"000000000000" when X = 290 AND Y = 47 else
"000000000000" when X = 291 AND Y = 47 else
"000000000000" when X = 292 AND Y = 47 else
"000000000000" when X = 293 AND Y = 47 else
"000000000000" when X = 294 AND Y = 47 else
"000000000000" when X = 295 AND Y = 47 else
"000000000000" when X = 296 AND Y = 47 else
"000000000000" when X = 297 AND Y = 47 else
"000000000000" when X = 298 AND Y = 47 else
"000000000000" when X = 299 AND Y = 47 else
"000000000000" when X = 300 AND Y = 47 else
"000000000000" when X = 301 AND Y = 47 else
"000000000000" when X = 302 AND Y = 47 else
"000000000000" when X = 303 AND Y = 47 else
"000000000000" when X = 304 AND Y = 47 else
"000000000000" when X = 305 AND Y = 47 else
"000000000000" when X = 306 AND Y = 47 else
"000000000000" when X = 307 AND Y = 47 else
"000000000000" when X = 308 AND Y = 47 else
"000000000000" when X = 309 AND Y = 47 else
"000000000000" when X = 310 AND Y = 47 else
"000000000000" when X = 311 AND Y = 47 else
"000000000000" when X = 312 AND Y = 47 else
"000000000000" when X = 313 AND Y = 47 else
"000000000000" when X = 314 AND Y = 47 else
"000000000000" when X = 315 AND Y = 47 else
"000000000000" when X = 316 AND Y = 47 else
"000000000000" when X = 317 AND Y = 47 else
"000000000000" when X = 318 AND Y = 47 else
"000000000000" when X = 319 AND Y = 47 else
"000000000000" when X = 320 AND Y = 47 else
"000000000000" when X = 321 AND Y = 47 else
"000000000000" when X = 322 AND Y = 47 else
"000000000000" when X = 323 AND Y = 47 else
"000000000000" when X = 324 AND Y = 47 else
"000000000000" when X = 0 AND Y = 48 else
"000000000000" when X = 1 AND Y = 48 else
"000000000000" when X = 2 AND Y = 48 else
"000000000000" when X = 3 AND Y = 48 else
"000000000000" when X = 4 AND Y = 48 else
"000000000000" when X = 5 AND Y = 48 else
"000000000000" when X = 6 AND Y = 48 else
"000000000000" when X = 7 AND Y = 48 else
"000000000000" when X = 8 AND Y = 48 else
"000000000000" when X = 9 AND Y = 48 else
"000000000000" when X = 10 AND Y = 48 else
"000000000000" when X = 11 AND Y = 48 else
"000000000000" when X = 12 AND Y = 48 else
"000000000000" when X = 13 AND Y = 48 else
"000000000000" when X = 14 AND Y = 48 else
"000000000000" when X = 15 AND Y = 48 else
"000000000000" when X = 16 AND Y = 48 else
"000000000000" when X = 17 AND Y = 48 else
"000000000000" when X = 18 AND Y = 48 else
"000000000000" when X = 19 AND Y = 48 else
"000000000000" when X = 20 AND Y = 48 else
"000000000000" when X = 21 AND Y = 48 else
"000000000000" when X = 22 AND Y = 48 else
"000000000000" when X = 23 AND Y = 48 else
"000000000000" when X = 24 AND Y = 48 else
"000000000000" when X = 25 AND Y = 48 else
"000000000000" when X = 26 AND Y = 48 else
"000000000000" when X = 27 AND Y = 48 else
"000000000000" when X = 28 AND Y = 48 else
"000000000000" when X = 29 AND Y = 48 else
"000000000000" when X = 30 AND Y = 48 else
"000000000000" when X = 31 AND Y = 48 else
"000000000000" when X = 32 AND Y = 48 else
"000000000000" when X = 33 AND Y = 48 else
"000000000000" when X = 34 AND Y = 48 else
"000000000000" when X = 35 AND Y = 48 else
"000000000000" when X = 36 AND Y = 48 else
"000000000000" when X = 37 AND Y = 48 else
"000000000000" when X = 38 AND Y = 48 else
"000000000000" when X = 39 AND Y = 48 else
"100010011101" when X = 40 AND Y = 48 else
"100010011101" when X = 41 AND Y = 48 else
"100010011101" when X = 42 AND Y = 48 else
"100010011101" when X = 43 AND Y = 48 else
"100010011101" when X = 44 AND Y = 48 else
"100010011101" when X = 45 AND Y = 48 else
"100010011101" when X = 46 AND Y = 48 else
"100010011101" when X = 47 AND Y = 48 else
"100010011101" when X = 48 AND Y = 48 else
"100010011101" when X = 49 AND Y = 48 else
"110111011111" when X = 50 AND Y = 48 else
"110111011111" when X = 51 AND Y = 48 else
"110111011111" when X = 52 AND Y = 48 else
"110111011111" when X = 53 AND Y = 48 else
"110111011111" when X = 54 AND Y = 48 else
"110111011111" when X = 55 AND Y = 48 else
"110111011111" when X = 56 AND Y = 48 else
"110111011111" when X = 57 AND Y = 48 else
"110111011111" when X = 58 AND Y = 48 else
"110111011111" when X = 59 AND Y = 48 else
"111111111111" when X = 60 AND Y = 48 else
"111111111111" when X = 61 AND Y = 48 else
"111111111111" when X = 62 AND Y = 48 else
"111111111111" when X = 63 AND Y = 48 else
"111111111111" when X = 64 AND Y = 48 else
"111111111111" when X = 65 AND Y = 48 else
"111111111111" when X = 66 AND Y = 48 else
"111111111111" when X = 67 AND Y = 48 else
"111111111111" when X = 68 AND Y = 48 else
"111111111111" when X = 69 AND Y = 48 else
"111111111111" when X = 70 AND Y = 48 else
"111111111111" when X = 71 AND Y = 48 else
"111111111111" when X = 72 AND Y = 48 else
"111111111111" when X = 73 AND Y = 48 else
"111111111111" when X = 74 AND Y = 48 else
"111111111111" when X = 75 AND Y = 48 else
"111111111111" when X = 76 AND Y = 48 else
"111111111111" when X = 77 AND Y = 48 else
"111111111111" when X = 78 AND Y = 48 else
"111111111111" when X = 79 AND Y = 48 else
"111111111111" when X = 80 AND Y = 48 else
"111111111111" when X = 81 AND Y = 48 else
"111111111111" when X = 82 AND Y = 48 else
"111111111111" when X = 83 AND Y = 48 else
"111111111111" when X = 84 AND Y = 48 else
"111111111111" when X = 85 AND Y = 48 else
"111111111111" when X = 86 AND Y = 48 else
"111111111111" when X = 87 AND Y = 48 else
"111111111111" when X = 88 AND Y = 48 else
"111111111111" when X = 89 AND Y = 48 else
"111111111111" when X = 90 AND Y = 48 else
"111111111111" when X = 91 AND Y = 48 else
"111111111111" when X = 92 AND Y = 48 else
"111111111111" when X = 93 AND Y = 48 else
"111111111111" when X = 94 AND Y = 48 else
"111111111111" when X = 95 AND Y = 48 else
"111111111111" when X = 96 AND Y = 48 else
"111111111111" when X = 97 AND Y = 48 else
"111111111111" when X = 98 AND Y = 48 else
"111111111111" when X = 99 AND Y = 48 else
"111111111111" when X = 100 AND Y = 48 else
"111111111111" when X = 101 AND Y = 48 else
"111111111111" when X = 102 AND Y = 48 else
"111111111111" when X = 103 AND Y = 48 else
"111111111111" when X = 104 AND Y = 48 else
"111111111111" when X = 105 AND Y = 48 else
"111111111111" when X = 106 AND Y = 48 else
"111111111111" when X = 107 AND Y = 48 else
"111111111111" when X = 108 AND Y = 48 else
"111111111111" when X = 109 AND Y = 48 else
"111111111111" when X = 110 AND Y = 48 else
"111111111111" when X = 111 AND Y = 48 else
"111111111111" when X = 112 AND Y = 48 else
"111111111111" when X = 113 AND Y = 48 else
"111111111111" when X = 114 AND Y = 48 else
"111111111111" when X = 115 AND Y = 48 else
"111111111111" when X = 116 AND Y = 48 else
"111111111111" when X = 117 AND Y = 48 else
"111111111111" when X = 118 AND Y = 48 else
"111111111111" when X = 119 AND Y = 48 else
"111111111111" when X = 120 AND Y = 48 else
"111111111111" when X = 121 AND Y = 48 else
"111111111111" when X = 122 AND Y = 48 else
"111111111111" when X = 123 AND Y = 48 else
"111111111111" when X = 124 AND Y = 48 else
"111111111111" when X = 125 AND Y = 48 else
"111111111111" when X = 126 AND Y = 48 else
"111111111111" when X = 127 AND Y = 48 else
"111111111111" when X = 128 AND Y = 48 else
"111111111111" when X = 129 AND Y = 48 else
"111111111111" when X = 130 AND Y = 48 else
"111111111111" when X = 131 AND Y = 48 else
"111111111111" when X = 132 AND Y = 48 else
"111111111111" when X = 133 AND Y = 48 else
"111111111111" when X = 134 AND Y = 48 else
"111111111111" when X = 135 AND Y = 48 else
"111111111111" when X = 136 AND Y = 48 else
"111111111111" when X = 137 AND Y = 48 else
"111111111111" when X = 138 AND Y = 48 else
"111111111111" when X = 139 AND Y = 48 else
"111111111111" when X = 140 AND Y = 48 else
"111111111111" when X = 141 AND Y = 48 else
"111111111111" when X = 142 AND Y = 48 else
"111111111111" when X = 143 AND Y = 48 else
"111111111111" when X = 144 AND Y = 48 else
"111111111111" when X = 145 AND Y = 48 else
"111111111111" when X = 146 AND Y = 48 else
"111111111111" when X = 147 AND Y = 48 else
"111111111111" when X = 148 AND Y = 48 else
"111111111111" when X = 149 AND Y = 48 else
"111111111111" when X = 150 AND Y = 48 else
"111111111111" when X = 151 AND Y = 48 else
"111111111111" when X = 152 AND Y = 48 else
"111111111111" when X = 153 AND Y = 48 else
"111111111111" when X = 154 AND Y = 48 else
"111111111111" when X = 155 AND Y = 48 else
"111111111111" when X = 156 AND Y = 48 else
"111111111111" when X = 157 AND Y = 48 else
"111111111111" when X = 158 AND Y = 48 else
"111111111111" when X = 159 AND Y = 48 else
"111111111111" when X = 160 AND Y = 48 else
"111111111111" when X = 161 AND Y = 48 else
"111111111111" when X = 162 AND Y = 48 else
"111111111111" when X = 163 AND Y = 48 else
"111111111111" when X = 164 AND Y = 48 else
"111111111111" when X = 165 AND Y = 48 else
"111111111111" when X = 166 AND Y = 48 else
"111111111111" when X = 167 AND Y = 48 else
"111111111111" when X = 168 AND Y = 48 else
"111111111111" when X = 169 AND Y = 48 else
"111111111111" when X = 170 AND Y = 48 else
"111111111111" when X = 171 AND Y = 48 else
"111111111111" when X = 172 AND Y = 48 else
"111111111111" when X = 173 AND Y = 48 else
"111111111111" when X = 174 AND Y = 48 else
"111111111111" when X = 175 AND Y = 48 else
"111111111111" when X = 176 AND Y = 48 else
"111111111111" when X = 177 AND Y = 48 else
"111111111111" when X = 178 AND Y = 48 else
"111111111111" when X = 179 AND Y = 48 else
"111111111111" when X = 180 AND Y = 48 else
"111111111111" when X = 181 AND Y = 48 else
"111111111111" when X = 182 AND Y = 48 else
"111111111111" when X = 183 AND Y = 48 else
"111111111111" when X = 184 AND Y = 48 else
"111111111111" when X = 185 AND Y = 48 else
"111111111111" when X = 186 AND Y = 48 else
"111111111111" when X = 187 AND Y = 48 else
"111111111111" when X = 188 AND Y = 48 else
"111111111111" when X = 189 AND Y = 48 else
"111111111111" when X = 190 AND Y = 48 else
"111111111111" when X = 191 AND Y = 48 else
"111111111111" when X = 192 AND Y = 48 else
"111111111111" when X = 193 AND Y = 48 else
"111111111111" when X = 194 AND Y = 48 else
"111111111111" when X = 195 AND Y = 48 else
"111111111111" when X = 196 AND Y = 48 else
"111111111111" when X = 197 AND Y = 48 else
"111111111111" when X = 198 AND Y = 48 else
"111111111111" when X = 199 AND Y = 48 else
"111111111111" when X = 200 AND Y = 48 else
"111111111111" when X = 201 AND Y = 48 else
"111111111111" when X = 202 AND Y = 48 else
"111111111111" when X = 203 AND Y = 48 else
"111111111111" when X = 204 AND Y = 48 else
"111111111111" when X = 205 AND Y = 48 else
"111111111111" when X = 206 AND Y = 48 else
"111111111111" when X = 207 AND Y = 48 else
"111111111111" when X = 208 AND Y = 48 else
"111111111111" when X = 209 AND Y = 48 else
"111111111111" when X = 210 AND Y = 48 else
"111111111111" when X = 211 AND Y = 48 else
"111111111111" when X = 212 AND Y = 48 else
"111111111111" when X = 213 AND Y = 48 else
"111111111111" when X = 214 AND Y = 48 else
"111111111111" when X = 215 AND Y = 48 else
"111111111111" when X = 216 AND Y = 48 else
"111111111111" when X = 217 AND Y = 48 else
"111111111111" when X = 218 AND Y = 48 else
"111111111111" when X = 219 AND Y = 48 else
"111111111111" when X = 220 AND Y = 48 else
"111111111111" when X = 221 AND Y = 48 else
"111111111111" when X = 222 AND Y = 48 else
"111111111111" when X = 223 AND Y = 48 else
"111111111111" when X = 224 AND Y = 48 else
"111111111111" when X = 225 AND Y = 48 else
"111111111111" when X = 226 AND Y = 48 else
"111111111111" when X = 227 AND Y = 48 else
"111111111111" when X = 228 AND Y = 48 else
"111111111111" when X = 229 AND Y = 48 else
"111111111111" when X = 230 AND Y = 48 else
"111111111111" when X = 231 AND Y = 48 else
"111111111111" when X = 232 AND Y = 48 else
"111111111111" when X = 233 AND Y = 48 else
"111111111111" when X = 234 AND Y = 48 else
"111111111111" when X = 235 AND Y = 48 else
"111111111111" when X = 236 AND Y = 48 else
"111111111111" when X = 237 AND Y = 48 else
"111111111111" when X = 238 AND Y = 48 else
"111111111111" when X = 239 AND Y = 48 else
"111111111111" when X = 240 AND Y = 48 else
"111111111111" when X = 241 AND Y = 48 else
"111111111111" when X = 242 AND Y = 48 else
"111111111111" when X = 243 AND Y = 48 else
"111111111111" when X = 244 AND Y = 48 else
"111111111111" when X = 245 AND Y = 48 else
"111111111111" when X = 246 AND Y = 48 else
"111111111111" when X = 247 AND Y = 48 else
"111111111111" when X = 248 AND Y = 48 else
"111111111111" when X = 249 AND Y = 48 else
"111111111111" when X = 250 AND Y = 48 else
"111111111111" when X = 251 AND Y = 48 else
"111111111111" when X = 252 AND Y = 48 else
"111111111111" when X = 253 AND Y = 48 else
"111111111111" when X = 254 AND Y = 48 else
"111111111111" when X = 255 AND Y = 48 else
"111111111111" when X = 256 AND Y = 48 else
"111111111111" when X = 257 AND Y = 48 else
"111111111111" when X = 258 AND Y = 48 else
"111111111111" when X = 259 AND Y = 48 else
"111111111111" when X = 260 AND Y = 48 else
"111111111111" when X = 261 AND Y = 48 else
"111111111111" when X = 262 AND Y = 48 else
"111111111111" when X = 263 AND Y = 48 else
"111111111111" when X = 264 AND Y = 48 else
"110111011111" when X = 265 AND Y = 48 else
"110111011111" when X = 266 AND Y = 48 else
"110111011111" when X = 267 AND Y = 48 else
"110111011111" when X = 268 AND Y = 48 else
"110111011111" when X = 269 AND Y = 48 else
"110111011111" when X = 270 AND Y = 48 else
"110111011111" when X = 271 AND Y = 48 else
"110111011111" when X = 272 AND Y = 48 else
"110111011111" when X = 273 AND Y = 48 else
"110111011111" when X = 274 AND Y = 48 else
"110111011111" when X = 275 AND Y = 48 else
"110111011111" when X = 276 AND Y = 48 else
"110111011111" when X = 277 AND Y = 48 else
"110111011111" when X = 278 AND Y = 48 else
"110111011111" when X = 279 AND Y = 48 else
"000000000000" when X = 280 AND Y = 48 else
"000000000000" when X = 281 AND Y = 48 else
"000000000000" when X = 282 AND Y = 48 else
"000000000000" when X = 283 AND Y = 48 else
"000000000000" when X = 284 AND Y = 48 else
"000000000000" when X = 285 AND Y = 48 else
"000000000000" when X = 286 AND Y = 48 else
"000000000000" when X = 287 AND Y = 48 else
"000000000000" when X = 288 AND Y = 48 else
"000000000000" when X = 289 AND Y = 48 else
"000000000000" when X = 290 AND Y = 48 else
"000000000000" when X = 291 AND Y = 48 else
"000000000000" when X = 292 AND Y = 48 else
"000000000000" when X = 293 AND Y = 48 else
"000000000000" when X = 294 AND Y = 48 else
"000000000000" when X = 295 AND Y = 48 else
"000000000000" when X = 296 AND Y = 48 else
"000000000000" when X = 297 AND Y = 48 else
"000000000000" when X = 298 AND Y = 48 else
"000000000000" when X = 299 AND Y = 48 else
"000000000000" when X = 300 AND Y = 48 else
"000000000000" when X = 301 AND Y = 48 else
"000000000000" when X = 302 AND Y = 48 else
"000000000000" when X = 303 AND Y = 48 else
"000000000000" when X = 304 AND Y = 48 else
"000000000000" when X = 305 AND Y = 48 else
"000000000000" when X = 306 AND Y = 48 else
"000000000000" when X = 307 AND Y = 48 else
"000000000000" when X = 308 AND Y = 48 else
"000000000000" when X = 309 AND Y = 48 else
"000000000000" when X = 310 AND Y = 48 else
"000000000000" when X = 311 AND Y = 48 else
"000000000000" when X = 312 AND Y = 48 else
"000000000000" when X = 313 AND Y = 48 else
"000000000000" when X = 314 AND Y = 48 else
"000000000000" when X = 315 AND Y = 48 else
"000000000000" when X = 316 AND Y = 48 else
"000000000000" when X = 317 AND Y = 48 else
"000000000000" when X = 318 AND Y = 48 else
"000000000000" when X = 319 AND Y = 48 else
"000000000000" when X = 320 AND Y = 48 else
"000000000000" when X = 321 AND Y = 48 else
"000000000000" when X = 322 AND Y = 48 else
"000000000000" when X = 323 AND Y = 48 else
"000000000000" when X = 324 AND Y = 48 else
"000000000000" when X = 0 AND Y = 49 else
"000000000000" when X = 1 AND Y = 49 else
"000000000000" when X = 2 AND Y = 49 else
"000000000000" when X = 3 AND Y = 49 else
"000000000000" when X = 4 AND Y = 49 else
"000000000000" when X = 5 AND Y = 49 else
"000000000000" when X = 6 AND Y = 49 else
"000000000000" when X = 7 AND Y = 49 else
"000000000000" when X = 8 AND Y = 49 else
"000000000000" when X = 9 AND Y = 49 else
"000000000000" when X = 10 AND Y = 49 else
"000000000000" when X = 11 AND Y = 49 else
"000000000000" when X = 12 AND Y = 49 else
"000000000000" when X = 13 AND Y = 49 else
"000000000000" when X = 14 AND Y = 49 else
"000000000000" when X = 15 AND Y = 49 else
"000000000000" when X = 16 AND Y = 49 else
"000000000000" when X = 17 AND Y = 49 else
"000000000000" when X = 18 AND Y = 49 else
"000000000000" when X = 19 AND Y = 49 else
"000000000000" when X = 20 AND Y = 49 else
"000000000000" when X = 21 AND Y = 49 else
"000000000000" when X = 22 AND Y = 49 else
"000000000000" when X = 23 AND Y = 49 else
"000000000000" when X = 24 AND Y = 49 else
"000000000000" when X = 25 AND Y = 49 else
"000000000000" when X = 26 AND Y = 49 else
"000000000000" when X = 27 AND Y = 49 else
"000000000000" when X = 28 AND Y = 49 else
"000000000000" when X = 29 AND Y = 49 else
"000000000000" when X = 30 AND Y = 49 else
"000000000000" when X = 31 AND Y = 49 else
"000000000000" when X = 32 AND Y = 49 else
"000000000000" when X = 33 AND Y = 49 else
"000000000000" when X = 34 AND Y = 49 else
"000000000000" when X = 35 AND Y = 49 else
"000000000000" when X = 36 AND Y = 49 else
"000000000000" when X = 37 AND Y = 49 else
"000000000000" when X = 38 AND Y = 49 else
"000000000000" when X = 39 AND Y = 49 else
"100010011101" when X = 40 AND Y = 49 else
"100010011101" when X = 41 AND Y = 49 else
"100010011101" when X = 42 AND Y = 49 else
"100010011101" when X = 43 AND Y = 49 else
"100010011101" when X = 44 AND Y = 49 else
"100010011101" when X = 45 AND Y = 49 else
"100010011101" when X = 46 AND Y = 49 else
"100010011101" when X = 47 AND Y = 49 else
"100010011101" when X = 48 AND Y = 49 else
"100010011101" when X = 49 AND Y = 49 else
"110111011111" when X = 50 AND Y = 49 else
"110111011111" when X = 51 AND Y = 49 else
"110111011111" when X = 52 AND Y = 49 else
"110111011111" when X = 53 AND Y = 49 else
"110111011111" when X = 54 AND Y = 49 else
"110111011111" when X = 55 AND Y = 49 else
"110111011111" when X = 56 AND Y = 49 else
"110111011111" when X = 57 AND Y = 49 else
"110111011111" when X = 58 AND Y = 49 else
"110111011111" when X = 59 AND Y = 49 else
"111111111111" when X = 60 AND Y = 49 else
"111111111111" when X = 61 AND Y = 49 else
"111111111111" when X = 62 AND Y = 49 else
"111111111111" when X = 63 AND Y = 49 else
"111111111111" when X = 64 AND Y = 49 else
"111111111111" when X = 65 AND Y = 49 else
"111111111111" when X = 66 AND Y = 49 else
"111111111111" when X = 67 AND Y = 49 else
"111111111111" when X = 68 AND Y = 49 else
"111111111111" when X = 69 AND Y = 49 else
"111111111111" when X = 70 AND Y = 49 else
"111111111111" when X = 71 AND Y = 49 else
"111111111111" when X = 72 AND Y = 49 else
"111111111111" when X = 73 AND Y = 49 else
"111111111111" when X = 74 AND Y = 49 else
"111111111111" when X = 75 AND Y = 49 else
"111111111111" when X = 76 AND Y = 49 else
"111111111111" when X = 77 AND Y = 49 else
"111111111111" when X = 78 AND Y = 49 else
"111111111111" when X = 79 AND Y = 49 else
"111111111111" when X = 80 AND Y = 49 else
"111111111111" when X = 81 AND Y = 49 else
"111111111111" when X = 82 AND Y = 49 else
"111111111111" when X = 83 AND Y = 49 else
"111111111111" when X = 84 AND Y = 49 else
"111111111111" when X = 85 AND Y = 49 else
"111111111111" when X = 86 AND Y = 49 else
"111111111111" when X = 87 AND Y = 49 else
"111111111111" when X = 88 AND Y = 49 else
"111111111111" when X = 89 AND Y = 49 else
"111111111111" when X = 90 AND Y = 49 else
"111111111111" when X = 91 AND Y = 49 else
"111111111111" when X = 92 AND Y = 49 else
"111111111111" when X = 93 AND Y = 49 else
"111111111111" when X = 94 AND Y = 49 else
"111111111111" when X = 95 AND Y = 49 else
"111111111111" when X = 96 AND Y = 49 else
"111111111111" when X = 97 AND Y = 49 else
"111111111111" when X = 98 AND Y = 49 else
"111111111111" when X = 99 AND Y = 49 else
"111111111111" when X = 100 AND Y = 49 else
"111111111111" when X = 101 AND Y = 49 else
"111111111111" when X = 102 AND Y = 49 else
"111111111111" when X = 103 AND Y = 49 else
"111111111111" when X = 104 AND Y = 49 else
"111111111111" when X = 105 AND Y = 49 else
"111111111111" when X = 106 AND Y = 49 else
"111111111111" when X = 107 AND Y = 49 else
"111111111111" when X = 108 AND Y = 49 else
"111111111111" when X = 109 AND Y = 49 else
"111111111111" when X = 110 AND Y = 49 else
"111111111111" when X = 111 AND Y = 49 else
"111111111111" when X = 112 AND Y = 49 else
"111111111111" when X = 113 AND Y = 49 else
"111111111111" when X = 114 AND Y = 49 else
"111111111111" when X = 115 AND Y = 49 else
"111111111111" when X = 116 AND Y = 49 else
"111111111111" when X = 117 AND Y = 49 else
"111111111111" when X = 118 AND Y = 49 else
"111111111111" when X = 119 AND Y = 49 else
"111111111111" when X = 120 AND Y = 49 else
"111111111111" when X = 121 AND Y = 49 else
"111111111111" when X = 122 AND Y = 49 else
"111111111111" when X = 123 AND Y = 49 else
"111111111111" when X = 124 AND Y = 49 else
"111111111111" when X = 125 AND Y = 49 else
"111111111111" when X = 126 AND Y = 49 else
"111111111111" when X = 127 AND Y = 49 else
"111111111111" when X = 128 AND Y = 49 else
"111111111111" when X = 129 AND Y = 49 else
"111111111111" when X = 130 AND Y = 49 else
"111111111111" when X = 131 AND Y = 49 else
"111111111111" when X = 132 AND Y = 49 else
"111111111111" when X = 133 AND Y = 49 else
"111111111111" when X = 134 AND Y = 49 else
"111111111111" when X = 135 AND Y = 49 else
"111111111111" when X = 136 AND Y = 49 else
"111111111111" when X = 137 AND Y = 49 else
"111111111111" when X = 138 AND Y = 49 else
"111111111111" when X = 139 AND Y = 49 else
"111111111111" when X = 140 AND Y = 49 else
"111111111111" when X = 141 AND Y = 49 else
"111111111111" when X = 142 AND Y = 49 else
"111111111111" when X = 143 AND Y = 49 else
"111111111111" when X = 144 AND Y = 49 else
"111111111111" when X = 145 AND Y = 49 else
"111111111111" when X = 146 AND Y = 49 else
"111111111111" when X = 147 AND Y = 49 else
"111111111111" when X = 148 AND Y = 49 else
"111111111111" when X = 149 AND Y = 49 else
"111111111111" when X = 150 AND Y = 49 else
"111111111111" when X = 151 AND Y = 49 else
"111111111111" when X = 152 AND Y = 49 else
"111111111111" when X = 153 AND Y = 49 else
"111111111111" when X = 154 AND Y = 49 else
"111111111111" when X = 155 AND Y = 49 else
"111111111111" when X = 156 AND Y = 49 else
"111111111111" when X = 157 AND Y = 49 else
"111111111111" when X = 158 AND Y = 49 else
"111111111111" when X = 159 AND Y = 49 else
"111111111111" when X = 160 AND Y = 49 else
"111111111111" when X = 161 AND Y = 49 else
"111111111111" when X = 162 AND Y = 49 else
"111111111111" when X = 163 AND Y = 49 else
"111111111111" when X = 164 AND Y = 49 else
"111111111111" when X = 165 AND Y = 49 else
"111111111111" when X = 166 AND Y = 49 else
"111111111111" when X = 167 AND Y = 49 else
"111111111111" when X = 168 AND Y = 49 else
"111111111111" when X = 169 AND Y = 49 else
"111111111111" when X = 170 AND Y = 49 else
"111111111111" when X = 171 AND Y = 49 else
"111111111111" when X = 172 AND Y = 49 else
"111111111111" when X = 173 AND Y = 49 else
"111111111111" when X = 174 AND Y = 49 else
"111111111111" when X = 175 AND Y = 49 else
"111111111111" when X = 176 AND Y = 49 else
"111111111111" when X = 177 AND Y = 49 else
"111111111111" when X = 178 AND Y = 49 else
"111111111111" when X = 179 AND Y = 49 else
"111111111111" when X = 180 AND Y = 49 else
"111111111111" when X = 181 AND Y = 49 else
"111111111111" when X = 182 AND Y = 49 else
"111111111111" when X = 183 AND Y = 49 else
"111111111111" when X = 184 AND Y = 49 else
"111111111111" when X = 185 AND Y = 49 else
"111111111111" when X = 186 AND Y = 49 else
"111111111111" when X = 187 AND Y = 49 else
"111111111111" when X = 188 AND Y = 49 else
"111111111111" when X = 189 AND Y = 49 else
"111111111111" when X = 190 AND Y = 49 else
"111111111111" when X = 191 AND Y = 49 else
"111111111111" when X = 192 AND Y = 49 else
"111111111111" when X = 193 AND Y = 49 else
"111111111111" when X = 194 AND Y = 49 else
"111111111111" when X = 195 AND Y = 49 else
"111111111111" when X = 196 AND Y = 49 else
"111111111111" when X = 197 AND Y = 49 else
"111111111111" when X = 198 AND Y = 49 else
"111111111111" when X = 199 AND Y = 49 else
"111111111111" when X = 200 AND Y = 49 else
"111111111111" when X = 201 AND Y = 49 else
"111111111111" when X = 202 AND Y = 49 else
"111111111111" when X = 203 AND Y = 49 else
"111111111111" when X = 204 AND Y = 49 else
"111111111111" when X = 205 AND Y = 49 else
"111111111111" when X = 206 AND Y = 49 else
"111111111111" when X = 207 AND Y = 49 else
"111111111111" when X = 208 AND Y = 49 else
"111111111111" when X = 209 AND Y = 49 else
"111111111111" when X = 210 AND Y = 49 else
"111111111111" when X = 211 AND Y = 49 else
"111111111111" when X = 212 AND Y = 49 else
"111111111111" when X = 213 AND Y = 49 else
"111111111111" when X = 214 AND Y = 49 else
"111111111111" when X = 215 AND Y = 49 else
"111111111111" when X = 216 AND Y = 49 else
"111111111111" when X = 217 AND Y = 49 else
"111111111111" when X = 218 AND Y = 49 else
"111111111111" when X = 219 AND Y = 49 else
"111111111111" when X = 220 AND Y = 49 else
"111111111111" when X = 221 AND Y = 49 else
"111111111111" when X = 222 AND Y = 49 else
"111111111111" when X = 223 AND Y = 49 else
"111111111111" when X = 224 AND Y = 49 else
"111111111111" when X = 225 AND Y = 49 else
"111111111111" when X = 226 AND Y = 49 else
"111111111111" when X = 227 AND Y = 49 else
"111111111111" when X = 228 AND Y = 49 else
"111111111111" when X = 229 AND Y = 49 else
"111111111111" when X = 230 AND Y = 49 else
"111111111111" when X = 231 AND Y = 49 else
"111111111111" when X = 232 AND Y = 49 else
"111111111111" when X = 233 AND Y = 49 else
"111111111111" when X = 234 AND Y = 49 else
"111111111111" when X = 235 AND Y = 49 else
"111111111111" when X = 236 AND Y = 49 else
"111111111111" when X = 237 AND Y = 49 else
"111111111111" when X = 238 AND Y = 49 else
"111111111111" when X = 239 AND Y = 49 else
"111111111111" when X = 240 AND Y = 49 else
"111111111111" when X = 241 AND Y = 49 else
"111111111111" when X = 242 AND Y = 49 else
"111111111111" when X = 243 AND Y = 49 else
"111111111111" when X = 244 AND Y = 49 else
"111111111111" when X = 245 AND Y = 49 else
"111111111111" when X = 246 AND Y = 49 else
"111111111111" when X = 247 AND Y = 49 else
"111111111111" when X = 248 AND Y = 49 else
"111111111111" when X = 249 AND Y = 49 else
"111111111111" when X = 250 AND Y = 49 else
"111111111111" when X = 251 AND Y = 49 else
"111111111111" when X = 252 AND Y = 49 else
"111111111111" when X = 253 AND Y = 49 else
"111111111111" when X = 254 AND Y = 49 else
"111111111111" when X = 255 AND Y = 49 else
"111111111111" when X = 256 AND Y = 49 else
"111111111111" when X = 257 AND Y = 49 else
"111111111111" when X = 258 AND Y = 49 else
"111111111111" when X = 259 AND Y = 49 else
"111111111111" when X = 260 AND Y = 49 else
"111111111111" when X = 261 AND Y = 49 else
"111111111111" when X = 262 AND Y = 49 else
"111111111111" when X = 263 AND Y = 49 else
"111111111111" when X = 264 AND Y = 49 else
"110111011111" when X = 265 AND Y = 49 else
"110111011111" when X = 266 AND Y = 49 else
"110111011111" when X = 267 AND Y = 49 else
"110111011111" when X = 268 AND Y = 49 else
"110111011111" when X = 269 AND Y = 49 else
"110111011111" when X = 270 AND Y = 49 else
"110111011111" when X = 271 AND Y = 49 else
"110111011111" when X = 272 AND Y = 49 else
"110111011111" when X = 273 AND Y = 49 else
"110111011111" when X = 274 AND Y = 49 else
"110111011111" when X = 275 AND Y = 49 else
"110111011111" when X = 276 AND Y = 49 else
"110111011111" when X = 277 AND Y = 49 else
"110111011111" when X = 278 AND Y = 49 else
"110111011111" when X = 279 AND Y = 49 else
"000000000000" when X = 280 AND Y = 49 else
"000000000000" when X = 281 AND Y = 49 else
"000000000000" when X = 282 AND Y = 49 else
"000000000000" when X = 283 AND Y = 49 else
"000000000000" when X = 284 AND Y = 49 else
"000000000000" when X = 285 AND Y = 49 else
"000000000000" when X = 286 AND Y = 49 else
"000000000000" when X = 287 AND Y = 49 else
"000000000000" when X = 288 AND Y = 49 else
"000000000000" when X = 289 AND Y = 49 else
"000000000000" when X = 290 AND Y = 49 else
"000000000000" when X = 291 AND Y = 49 else
"000000000000" when X = 292 AND Y = 49 else
"000000000000" when X = 293 AND Y = 49 else
"000000000000" when X = 294 AND Y = 49 else
"000000000000" when X = 295 AND Y = 49 else
"000000000000" when X = 296 AND Y = 49 else
"000000000000" when X = 297 AND Y = 49 else
"000000000000" when X = 298 AND Y = 49 else
"000000000000" when X = 299 AND Y = 49 else
"000000000000" when X = 300 AND Y = 49 else
"000000000000" when X = 301 AND Y = 49 else
"000000000000" when X = 302 AND Y = 49 else
"000000000000" when X = 303 AND Y = 49 else
"000000000000" when X = 304 AND Y = 49 else
"000000000000" when X = 305 AND Y = 49 else
"000000000000" when X = 306 AND Y = 49 else
"000000000000" when X = 307 AND Y = 49 else
"000000000000" when X = 308 AND Y = 49 else
"000000000000" when X = 309 AND Y = 49 else
"000000000000" when X = 310 AND Y = 49 else
"000000000000" when X = 311 AND Y = 49 else
"000000000000" when X = 312 AND Y = 49 else
"000000000000" when X = 313 AND Y = 49 else
"000000000000" when X = 314 AND Y = 49 else
"000000000000" when X = 315 AND Y = 49 else
"000000000000" when X = 316 AND Y = 49 else
"000000000000" when X = 317 AND Y = 49 else
"000000000000" when X = 318 AND Y = 49 else
"000000000000" when X = 319 AND Y = 49 else
"000000000000" when X = 320 AND Y = 49 else
"000000000000" when X = 321 AND Y = 49 else
"000000000000" when X = 322 AND Y = 49 else
"000000000000" when X = 323 AND Y = 49 else
"000000000000" when X = 324 AND Y = 49 else
"100010011101" when X = 0 AND Y = 50 else
"100010011101" when X = 1 AND Y = 50 else
"100010011101" when X = 2 AND Y = 50 else
"100010011101" when X = 3 AND Y = 50 else
"100010011101" when X = 4 AND Y = 50 else
"100010011101" when X = 5 AND Y = 50 else
"100010011101" when X = 6 AND Y = 50 else
"100010011101" when X = 7 AND Y = 50 else
"100010011101" when X = 8 AND Y = 50 else
"100010011101" when X = 9 AND Y = 50 else
"100010011101" when X = 10 AND Y = 50 else
"100010011101" when X = 11 AND Y = 50 else
"100010011101" when X = 12 AND Y = 50 else
"100010011101" when X = 13 AND Y = 50 else
"100010011101" when X = 14 AND Y = 50 else
"100010011101" when X = 15 AND Y = 50 else
"100010011101" when X = 16 AND Y = 50 else
"100010011101" when X = 17 AND Y = 50 else
"100010011101" when X = 18 AND Y = 50 else
"100010011101" when X = 19 AND Y = 50 else
"100010011101" when X = 20 AND Y = 50 else
"100010011101" when X = 21 AND Y = 50 else
"100010011101" when X = 22 AND Y = 50 else
"100010011101" when X = 23 AND Y = 50 else
"100010011101" when X = 24 AND Y = 50 else
"100010011101" when X = 25 AND Y = 50 else
"100010011101" when X = 26 AND Y = 50 else
"100010011101" when X = 27 AND Y = 50 else
"100010011101" when X = 28 AND Y = 50 else
"100010011101" when X = 29 AND Y = 50 else
"100010011101" when X = 30 AND Y = 50 else
"100010011101" when X = 31 AND Y = 50 else
"100010011101" when X = 32 AND Y = 50 else
"100010011101" when X = 33 AND Y = 50 else
"100010011101" when X = 34 AND Y = 50 else
"100010011101" when X = 35 AND Y = 50 else
"100010011101" when X = 36 AND Y = 50 else
"100010011101" when X = 37 AND Y = 50 else
"100010011101" when X = 38 AND Y = 50 else
"100010011101" when X = 39 AND Y = 50 else
"100010011101" when X = 40 AND Y = 50 else
"100010011101" when X = 41 AND Y = 50 else
"100010011101" when X = 42 AND Y = 50 else
"100010011101" when X = 43 AND Y = 50 else
"100010011101" when X = 44 AND Y = 50 else
"110111011111" when X = 45 AND Y = 50 else
"110111011111" when X = 46 AND Y = 50 else
"110111011111" when X = 47 AND Y = 50 else
"110111011111" when X = 48 AND Y = 50 else
"110111011111" when X = 49 AND Y = 50 else
"110111011111" when X = 50 AND Y = 50 else
"110111011111" when X = 51 AND Y = 50 else
"110111011111" when X = 52 AND Y = 50 else
"110111011111" when X = 53 AND Y = 50 else
"110111011111" when X = 54 AND Y = 50 else
"110111011111" when X = 55 AND Y = 50 else
"110111011111" when X = 56 AND Y = 50 else
"110111011111" when X = 57 AND Y = 50 else
"110111011111" when X = 58 AND Y = 50 else
"110111011111" when X = 59 AND Y = 50 else
"110111011111" when X = 60 AND Y = 50 else
"110111011111" when X = 61 AND Y = 50 else
"110111011111" when X = 62 AND Y = 50 else
"110111011111" when X = 63 AND Y = 50 else
"110111011111" when X = 64 AND Y = 50 else
"110111011111" when X = 65 AND Y = 50 else
"110111011111" when X = 66 AND Y = 50 else
"110111011111" when X = 67 AND Y = 50 else
"110111011111" when X = 68 AND Y = 50 else
"110111011111" when X = 69 AND Y = 50 else
"111111111111" when X = 70 AND Y = 50 else
"111111111111" when X = 71 AND Y = 50 else
"111111111111" when X = 72 AND Y = 50 else
"111111111111" when X = 73 AND Y = 50 else
"111111111111" when X = 74 AND Y = 50 else
"111111111111" when X = 75 AND Y = 50 else
"111111111111" when X = 76 AND Y = 50 else
"111111111111" when X = 77 AND Y = 50 else
"111111111111" when X = 78 AND Y = 50 else
"111111111111" when X = 79 AND Y = 50 else
"111111111111" when X = 80 AND Y = 50 else
"111111111111" when X = 81 AND Y = 50 else
"111111111111" when X = 82 AND Y = 50 else
"111111111111" when X = 83 AND Y = 50 else
"111111111111" when X = 84 AND Y = 50 else
"111111111111" when X = 85 AND Y = 50 else
"111111111111" when X = 86 AND Y = 50 else
"111111111111" when X = 87 AND Y = 50 else
"111111111111" when X = 88 AND Y = 50 else
"111111111111" when X = 89 AND Y = 50 else
"111111111111" when X = 90 AND Y = 50 else
"111111111111" when X = 91 AND Y = 50 else
"111111111111" when X = 92 AND Y = 50 else
"111111111111" when X = 93 AND Y = 50 else
"111111111111" when X = 94 AND Y = 50 else
"111111111111" when X = 95 AND Y = 50 else
"111111111111" when X = 96 AND Y = 50 else
"111111111111" when X = 97 AND Y = 50 else
"111111111111" when X = 98 AND Y = 50 else
"111111111111" when X = 99 AND Y = 50 else
"111111111111" when X = 100 AND Y = 50 else
"111111111111" when X = 101 AND Y = 50 else
"111111111111" when X = 102 AND Y = 50 else
"111111111111" when X = 103 AND Y = 50 else
"111111111111" when X = 104 AND Y = 50 else
"111111111111" when X = 105 AND Y = 50 else
"111111111111" when X = 106 AND Y = 50 else
"111111111111" when X = 107 AND Y = 50 else
"111111111111" when X = 108 AND Y = 50 else
"111111111111" when X = 109 AND Y = 50 else
"111111111111" when X = 110 AND Y = 50 else
"111111111111" when X = 111 AND Y = 50 else
"111111111111" when X = 112 AND Y = 50 else
"111111111111" when X = 113 AND Y = 50 else
"111111111111" when X = 114 AND Y = 50 else
"111111111111" when X = 115 AND Y = 50 else
"111111111111" when X = 116 AND Y = 50 else
"111111111111" when X = 117 AND Y = 50 else
"111111111111" when X = 118 AND Y = 50 else
"111111111111" when X = 119 AND Y = 50 else
"111111111111" when X = 120 AND Y = 50 else
"111111111111" when X = 121 AND Y = 50 else
"111111111111" when X = 122 AND Y = 50 else
"111111111111" when X = 123 AND Y = 50 else
"111111111111" when X = 124 AND Y = 50 else
"111111111111" when X = 125 AND Y = 50 else
"111111111111" when X = 126 AND Y = 50 else
"111111111111" when X = 127 AND Y = 50 else
"111111111111" when X = 128 AND Y = 50 else
"111111111111" when X = 129 AND Y = 50 else
"111111111111" when X = 130 AND Y = 50 else
"111111111111" when X = 131 AND Y = 50 else
"111111111111" when X = 132 AND Y = 50 else
"111111111111" when X = 133 AND Y = 50 else
"111111111111" when X = 134 AND Y = 50 else
"111111111111" when X = 135 AND Y = 50 else
"111111111111" when X = 136 AND Y = 50 else
"111111111111" when X = 137 AND Y = 50 else
"111111111111" when X = 138 AND Y = 50 else
"111111111111" when X = 139 AND Y = 50 else
"111111111111" when X = 140 AND Y = 50 else
"111111111111" when X = 141 AND Y = 50 else
"111111111111" when X = 142 AND Y = 50 else
"111111111111" when X = 143 AND Y = 50 else
"111111111111" when X = 144 AND Y = 50 else
"111111111111" when X = 145 AND Y = 50 else
"111111111111" when X = 146 AND Y = 50 else
"111111111111" when X = 147 AND Y = 50 else
"111111111111" when X = 148 AND Y = 50 else
"111111111111" when X = 149 AND Y = 50 else
"111111111111" when X = 150 AND Y = 50 else
"111111111111" when X = 151 AND Y = 50 else
"111111111111" when X = 152 AND Y = 50 else
"111111111111" when X = 153 AND Y = 50 else
"111111111111" when X = 154 AND Y = 50 else
"111111111111" when X = 155 AND Y = 50 else
"111111111111" when X = 156 AND Y = 50 else
"111111111111" when X = 157 AND Y = 50 else
"111111111111" when X = 158 AND Y = 50 else
"111111111111" when X = 159 AND Y = 50 else
"111111111111" when X = 160 AND Y = 50 else
"111111111111" when X = 161 AND Y = 50 else
"111111111111" when X = 162 AND Y = 50 else
"111111111111" when X = 163 AND Y = 50 else
"111111111111" when X = 164 AND Y = 50 else
"111111111111" when X = 165 AND Y = 50 else
"111111111111" when X = 166 AND Y = 50 else
"111111111111" when X = 167 AND Y = 50 else
"111111111111" when X = 168 AND Y = 50 else
"111111111111" when X = 169 AND Y = 50 else
"111111111111" when X = 170 AND Y = 50 else
"111111111111" when X = 171 AND Y = 50 else
"111111111111" when X = 172 AND Y = 50 else
"111111111111" when X = 173 AND Y = 50 else
"111111111111" when X = 174 AND Y = 50 else
"111111111111" when X = 175 AND Y = 50 else
"111111111111" when X = 176 AND Y = 50 else
"111111111111" when X = 177 AND Y = 50 else
"111111111111" when X = 178 AND Y = 50 else
"111111111111" when X = 179 AND Y = 50 else
"111111111111" when X = 180 AND Y = 50 else
"111111111111" when X = 181 AND Y = 50 else
"111111111111" when X = 182 AND Y = 50 else
"111111111111" when X = 183 AND Y = 50 else
"111111111111" when X = 184 AND Y = 50 else
"111111111111" when X = 185 AND Y = 50 else
"111111111111" when X = 186 AND Y = 50 else
"111111111111" when X = 187 AND Y = 50 else
"111111111111" when X = 188 AND Y = 50 else
"111111111111" when X = 189 AND Y = 50 else
"111111111111" when X = 190 AND Y = 50 else
"111111111111" when X = 191 AND Y = 50 else
"111111111111" when X = 192 AND Y = 50 else
"111111111111" when X = 193 AND Y = 50 else
"111111111111" when X = 194 AND Y = 50 else
"111111111111" when X = 195 AND Y = 50 else
"111111111111" when X = 196 AND Y = 50 else
"111111111111" when X = 197 AND Y = 50 else
"111111111111" when X = 198 AND Y = 50 else
"111111111111" when X = 199 AND Y = 50 else
"111111111111" when X = 200 AND Y = 50 else
"111111111111" when X = 201 AND Y = 50 else
"111111111111" when X = 202 AND Y = 50 else
"111111111111" when X = 203 AND Y = 50 else
"111111111111" when X = 204 AND Y = 50 else
"111111111111" when X = 205 AND Y = 50 else
"111111111111" when X = 206 AND Y = 50 else
"111111111111" when X = 207 AND Y = 50 else
"111111111111" when X = 208 AND Y = 50 else
"111111111111" when X = 209 AND Y = 50 else
"111111111111" when X = 210 AND Y = 50 else
"111111111111" when X = 211 AND Y = 50 else
"111111111111" when X = 212 AND Y = 50 else
"111111111111" when X = 213 AND Y = 50 else
"111111111111" when X = 214 AND Y = 50 else
"111111111111" when X = 215 AND Y = 50 else
"111111111111" when X = 216 AND Y = 50 else
"111111111111" when X = 217 AND Y = 50 else
"111111111111" when X = 218 AND Y = 50 else
"111111111111" when X = 219 AND Y = 50 else
"111111111111" when X = 220 AND Y = 50 else
"111111111111" when X = 221 AND Y = 50 else
"111111111111" when X = 222 AND Y = 50 else
"111111111111" when X = 223 AND Y = 50 else
"111111111111" when X = 224 AND Y = 50 else
"111111111111" when X = 225 AND Y = 50 else
"111111111111" when X = 226 AND Y = 50 else
"111111111111" when X = 227 AND Y = 50 else
"111111111111" when X = 228 AND Y = 50 else
"111111111111" when X = 229 AND Y = 50 else
"111111111111" when X = 230 AND Y = 50 else
"111111111111" when X = 231 AND Y = 50 else
"111111111111" when X = 232 AND Y = 50 else
"111111111111" when X = 233 AND Y = 50 else
"111111111111" when X = 234 AND Y = 50 else
"111111111111" when X = 235 AND Y = 50 else
"111111111111" when X = 236 AND Y = 50 else
"111111111111" when X = 237 AND Y = 50 else
"111111111111" when X = 238 AND Y = 50 else
"111111111111" when X = 239 AND Y = 50 else
"111111111111" when X = 240 AND Y = 50 else
"111111111111" when X = 241 AND Y = 50 else
"111111111111" when X = 242 AND Y = 50 else
"111111111111" when X = 243 AND Y = 50 else
"111111111111" when X = 244 AND Y = 50 else
"111111111111" when X = 245 AND Y = 50 else
"111111111111" when X = 246 AND Y = 50 else
"111111111111" when X = 247 AND Y = 50 else
"111111111111" when X = 248 AND Y = 50 else
"111111111111" when X = 249 AND Y = 50 else
"111111111111" when X = 250 AND Y = 50 else
"111111111111" when X = 251 AND Y = 50 else
"111111111111" when X = 252 AND Y = 50 else
"111111111111" when X = 253 AND Y = 50 else
"111111111111" when X = 254 AND Y = 50 else
"111111111111" when X = 255 AND Y = 50 else
"111111111111" when X = 256 AND Y = 50 else
"111111111111" when X = 257 AND Y = 50 else
"111111111111" when X = 258 AND Y = 50 else
"111111111111" when X = 259 AND Y = 50 else
"111111111111" when X = 260 AND Y = 50 else
"111111111111" when X = 261 AND Y = 50 else
"111111111111" when X = 262 AND Y = 50 else
"111111111111" when X = 263 AND Y = 50 else
"111111111111" when X = 264 AND Y = 50 else
"110111011111" when X = 265 AND Y = 50 else
"110111011111" when X = 266 AND Y = 50 else
"110111011111" when X = 267 AND Y = 50 else
"110111011111" when X = 268 AND Y = 50 else
"110111011111" when X = 269 AND Y = 50 else
"110111011111" when X = 270 AND Y = 50 else
"110111011111" when X = 271 AND Y = 50 else
"110111011111" when X = 272 AND Y = 50 else
"110111011111" when X = 273 AND Y = 50 else
"110111011111" when X = 274 AND Y = 50 else
"110111011111" when X = 275 AND Y = 50 else
"110111011111" when X = 276 AND Y = 50 else
"110111011111" when X = 277 AND Y = 50 else
"110111011111" when X = 278 AND Y = 50 else
"110111011111" when X = 279 AND Y = 50 else
"000000000000" when X = 280 AND Y = 50 else
"000000000000" when X = 281 AND Y = 50 else
"000000000000" when X = 282 AND Y = 50 else
"000000000000" when X = 283 AND Y = 50 else
"000000000000" when X = 284 AND Y = 50 else
"000000000000" when X = 285 AND Y = 50 else
"000000000000" when X = 286 AND Y = 50 else
"000000000000" when X = 287 AND Y = 50 else
"000000000000" when X = 288 AND Y = 50 else
"000000000000" when X = 289 AND Y = 50 else
"000000000000" when X = 290 AND Y = 50 else
"000000000000" when X = 291 AND Y = 50 else
"000000000000" when X = 292 AND Y = 50 else
"000000000000" when X = 293 AND Y = 50 else
"000000000000" when X = 294 AND Y = 50 else
"000000000000" when X = 295 AND Y = 50 else
"000000000000" when X = 296 AND Y = 50 else
"000000000000" when X = 297 AND Y = 50 else
"000000000000" when X = 298 AND Y = 50 else
"000000000000" when X = 299 AND Y = 50 else
"000000000000" when X = 300 AND Y = 50 else
"000000000000" when X = 301 AND Y = 50 else
"000000000000" when X = 302 AND Y = 50 else
"000000000000" when X = 303 AND Y = 50 else
"000000000000" when X = 304 AND Y = 50 else
"000000000000" when X = 305 AND Y = 50 else
"000000000000" when X = 306 AND Y = 50 else
"000000000000" when X = 307 AND Y = 50 else
"000000000000" when X = 308 AND Y = 50 else
"000000000000" when X = 309 AND Y = 50 else
"000000000000" when X = 310 AND Y = 50 else
"000000000000" when X = 311 AND Y = 50 else
"000000000000" when X = 312 AND Y = 50 else
"000000000000" when X = 313 AND Y = 50 else
"000000000000" when X = 314 AND Y = 50 else
"000000000000" when X = 315 AND Y = 50 else
"000000000000" when X = 316 AND Y = 50 else
"000000000000" when X = 317 AND Y = 50 else
"000000000000" when X = 318 AND Y = 50 else
"000000000000" when X = 319 AND Y = 50 else
"000000000000" when X = 320 AND Y = 50 else
"000000000000" when X = 321 AND Y = 50 else
"000000000000" when X = 322 AND Y = 50 else
"000000000000" when X = 323 AND Y = 50 else
"000000000000" when X = 324 AND Y = 50 else
"100010011101" when X = 0 AND Y = 51 else
"100010011101" when X = 1 AND Y = 51 else
"100010011101" when X = 2 AND Y = 51 else
"100010011101" when X = 3 AND Y = 51 else
"100010011101" when X = 4 AND Y = 51 else
"100010011101" when X = 5 AND Y = 51 else
"100010011101" when X = 6 AND Y = 51 else
"100010011101" when X = 7 AND Y = 51 else
"100010011101" when X = 8 AND Y = 51 else
"100010011101" when X = 9 AND Y = 51 else
"100010011101" when X = 10 AND Y = 51 else
"100010011101" when X = 11 AND Y = 51 else
"100010011101" when X = 12 AND Y = 51 else
"100010011101" when X = 13 AND Y = 51 else
"100010011101" when X = 14 AND Y = 51 else
"100010011101" when X = 15 AND Y = 51 else
"100010011101" when X = 16 AND Y = 51 else
"100010011101" when X = 17 AND Y = 51 else
"100010011101" when X = 18 AND Y = 51 else
"100010011101" when X = 19 AND Y = 51 else
"100010011101" when X = 20 AND Y = 51 else
"100010011101" when X = 21 AND Y = 51 else
"100010011101" when X = 22 AND Y = 51 else
"100010011101" when X = 23 AND Y = 51 else
"100010011101" when X = 24 AND Y = 51 else
"100010011101" when X = 25 AND Y = 51 else
"100010011101" when X = 26 AND Y = 51 else
"100010011101" when X = 27 AND Y = 51 else
"100010011101" when X = 28 AND Y = 51 else
"100010011101" when X = 29 AND Y = 51 else
"100010011101" when X = 30 AND Y = 51 else
"100010011101" when X = 31 AND Y = 51 else
"100010011101" when X = 32 AND Y = 51 else
"100010011101" when X = 33 AND Y = 51 else
"100010011101" when X = 34 AND Y = 51 else
"100010011101" when X = 35 AND Y = 51 else
"100010011101" when X = 36 AND Y = 51 else
"100010011101" when X = 37 AND Y = 51 else
"100010011101" when X = 38 AND Y = 51 else
"100010011101" when X = 39 AND Y = 51 else
"100010011101" when X = 40 AND Y = 51 else
"100010011101" when X = 41 AND Y = 51 else
"100010011101" when X = 42 AND Y = 51 else
"100010011101" when X = 43 AND Y = 51 else
"100010011101" when X = 44 AND Y = 51 else
"110111011111" when X = 45 AND Y = 51 else
"110111011111" when X = 46 AND Y = 51 else
"110111011111" when X = 47 AND Y = 51 else
"110111011111" when X = 48 AND Y = 51 else
"110111011111" when X = 49 AND Y = 51 else
"110111011111" when X = 50 AND Y = 51 else
"110111011111" when X = 51 AND Y = 51 else
"110111011111" when X = 52 AND Y = 51 else
"110111011111" when X = 53 AND Y = 51 else
"110111011111" when X = 54 AND Y = 51 else
"110111011111" when X = 55 AND Y = 51 else
"110111011111" when X = 56 AND Y = 51 else
"110111011111" when X = 57 AND Y = 51 else
"110111011111" when X = 58 AND Y = 51 else
"110111011111" when X = 59 AND Y = 51 else
"110111011111" when X = 60 AND Y = 51 else
"110111011111" when X = 61 AND Y = 51 else
"110111011111" when X = 62 AND Y = 51 else
"110111011111" when X = 63 AND Y = 51 else
"110111011111" when X = 64 AND Y = 51 else
"110111011111" when X = 65 AND Y = 51 else
"110111011111" when X = 66 AND Y = 51 else
"110111011111" when X = 67 AND Y = 51 else
"110111011111" when X = 68 AND Y = 51 else
"110111011111" when X = 69 AND Y = 51 else
"111111111111" when X = 70 AND Y = 51 else
"111111111111" when X = 71 AND Y = 51 else
"111111111111" when X = 72 AND Y = 51 else
"111111111111" when X = 73 AND Y = 51 else
"111111111111" when X = 74 AND Y = 51 else
"111111111111" when X = 75 AND Y = 51 else
"111111111111" when X = 76 AND Y = 51 else
"111111111111" when X = 77 AND Y = 51 else
"111111111111" when X = 78 AND Y = 51 else
"111111111111" when X = 79 AND Y = 51 else
"111111111111" when X = 80 AND Y = 51 else
"111111111111" when X = 81 AND Y = 51 else
"111111111111" when X = 82 AND Y = 51 else
"111111111111" when X = 83 AND Y = 51 else
"111111111111" when X = 84 AND Y = 51 else
"111111111111" when X = 85 AND Y = 51 else
"111111111111" when X = 86 AND Y = 51 else
"111111111111" when X = 87 AND Y = 51 else
"111111111111" when X = 88 AND Y = 51 else
"111111111111" when X = 89 AND Y = 51 else
"111111111111" when X = 90 AND Y = 51 else
"111111111111" when X = 91 AND Y = 51 else
"111111111111" when X = 92 AND Y = 51 else
"111111111111" when X = 93 AND Y = 51 else
"111111111111" when X = 94 AND Y = 51 else
"111111111111" when X = 95 AND Y = 51 else
"111111111111" when X = 96 AND Y = 51 else
"111111111111" when X = 97 AND Y = 51 else
"111111111111" when X = 98 AND Y = 51 else
"111111111111" when X = 99 AND Y = 51 else
"111111111111" when X = 100 AND Y = 51 else
"111111111111" when X = 101 AND Y = 51 else
"111111111111" when X = 102 AND Y = 51 else
"111111111111" when X = 103 AND Y = 51 else
"111111111111" when X = 104 AND Y = 51 else
"111111111111" when X = 105 AND Y = 51 else
"111111111111" when X = 106 AND Y = 51 else
"111111111111" when X = 107 AND Y = 51 else
"111111111111" when X = 108 AND Y = 51 else
"111111111111" when X = 109 AND Y = 51 else
"111111111111" when X = 110 AND Y = 51 else
"111111111111" when X = 111 AND Y = 51 else
"111111111111" when X = 112 AND Y = 51 else
"111111111111" when X = 113 AND Y = 51 else
"111111111111" when X = 114 AND Y = 51 else
"111111111111" when X = 115 AND Y = 51 else
"111111111111" when X = 116 AND Y = 51 else
"111111111111" when X = 117 AND Y = 51 else
"111111111111" when X = 118 AND Y = 51 else
"111111111111" when X = 119 AND Y = 51 else
"111111111111" when X = 120 AND Y = 51 else
"111111111111" when X = 121 AND Y = 51 else
"111111111111" when X = 122 AND Y = 51 else
"111111111111" when X = 123 AND Y = 51 else
"111111111111" when X = 124 AND Y = 51 else
"111111111111" when X = 125 AND Y = 51 else
"111111111111" when X = 126 AND Y = 51 else
"111111111111" when X = 127 AND Y = 51 else
"111111111111" when X = 128 AND Y = 51 else
"111111111111" when X = 129 AND Y = 51 else
"111111111111" when X = 130 AND Y = 51 else
"111111111111" when X = 131 AND Y = 51 else
"111111111111" when X = 132 AND Y = 51 else
"111111111111" when X = 133 AND Y = 51 else
"111111111111" when X = 134 AND Y = 51 else
"111111111111" when X = 135 AND Y = 51 else
"111111111111" when X = 136 AND Y = 51 else
"111111111111" when X = 137 AND Y = 51 else
"111111111111" when X = 138 AND Y = 51 else
"111111111111" when X = 139 AND Y = 51 else
"111111111111" when X = 140 AND Y = 51 else
"111111111111" when X = 141 AND Y = 51 else
"111111111111" when X = 142 AND Y = 51 else
"111111111111" when X = 143 AND Y = 51 else
"111111111111" when X = 144 AND Y = 51 else
"111111111111" when X = 145 AND Y = 51 else
"111111111111" when X = 146 AND Y = 51 else
"111111111111" when X = 147 AND Y = 51 else
"111111111111" when X = 148 AND Y = 51 else
"111111111111" when X = 149 AND Y = 51 else
"111111111111" when X = 150 AND Y = 51 else
"111111111111" when X = 151 AND Y = 51 else
"111111111111" when X = 152 AND Y = 51 else
"111111111111" when X = 153 AND Y = 51 else
"111111111111" when X = 154 AND Y = 51 else
"111111111111" when X = 155 AND Y = 51 else
"111111111111" when X = 156 AND Y = 51 else
"111111111111" when X = 157 AND Y = 51 else
"111111111111" when X = 158 AND Y = 51 else
"111111111111" when X = 159 AND Y = 51 else
"111111111111" when X = 160 AND Y = 51 else
"111111111111" when X = 161 AND Y = 51 else
"111111111111" when X = 162 AND Y = 51 else
"111111111111" when X = 163 AND Y = 51 else
"111111111111" when X = 164 AND Y = 51 else
"111111111111" when X = 165 AND Y = 51 else
"111111111111" when X = 166 AND Y = 51 else
"111111111111" when X = 167 AND Y = 51 else
"111111111111" when X = 168 AND Y = 51 else
"111111111111" when X = 169 AND Y = 51 else
"111111111111" when X = 170 AND Y = 51 else
"111111111111" when X = 171 AND Y = 51 else
"111111111111" when X = 172 AND Y = 51 else
"111111111111" when X = 173 AND Y = 51 else
"111111111111" when X = 174 AND Y = 51 else
"111111111111" when X = 175 AND Y = 51 else
"111111111111" when X = 176 AND Y = 51 else
"111111111111" when X = 177 AND Y = 51 else
"111111111111" when X = 178 AND Y = 51 else
"111111111111" when X = 179 AND Y = 51 else
"111111111111" when X = 180 AND Y = 51 else
"111111111111" when X = 181 AND Y = 51 else
"111111111111" when X = 182 AND Y = 51 else
"111111111111" when X = 183 AND Y = 51 else
"111111111111" when X = 184 AND Y = 51 else
"111111111111" when X = 185 AND Y = 51 else
"111111111111" when X = 186 AND Y = 51 else
"111111111111" when X = 187 AND Y = 51 else
"111111111111" when X = 188 AND Y = 51 else
"111111111111" when X = 189 AND Y = 51 else
"111111111111" when X = 190 AND Y = 51 else
"111111111111" when X = 191 AND Y = 51 else
"111111111111" when X = 192 AND Y = 51 else
"111111111111" when X = 193 AND Y = 51 else
"111111111111" when X = 194 AND Y = 51 else
"111111111111" when X = 195 AND Y = 51 else
"111111111111" when X = 196 AND Y = 51 else
"111111111111" when X = 197 AND Y = 51 else
"111111111111" when X = 198 AND Y = 51 else
"111111111111" when X = 199 AND Y = 51 else
"111111111111" when X = 200 AND Y = 51 else
"111111111111" when X = 201 AND Y = 51 else
"111111111111" when X = 202 AND Y = 51 else
"111111111111" when X = 203 AND Y = 51 else
"111111111111" when X = 204 AND Y = 51 else
"111111111111" when X = 205 AND Y = 51 else
"111111111111" when X = 206 AND Y = 51 else
"111111111111" when X = 207 AND Y = 51 else
"111111111111" when X = 208 AND Y = 51 else
"111111111111" when X = 209 AND Y = 51 else
"111111111111" when X = 210 AND Y = 51 else
"111111111111" when X = 211 AND Y = 51 else
"111111111111" when X = 212 AND Y = 51 else
"111111111111" when X = 213 AND Y = 51 else
"111111111111" when X = 214 AND Y = 51 else
"111111111111" when X = 215 AND Y = 51 else
"111111111111" when X = 216 AND Y = 51 else
"111111111111" when X = 217 AND Y = 51 else
"111111111111" when X = 218 AND Y = 51 else
"111111111111" when X = 219 AND Y = 51 else
"111111111111" when X = 220 AND Y = 51 else
"111111111111" when X = 221 AND Y = 51 else
"111111111111" when X = 222 AND Y = 51 else
"111111111111" when X = 223 AND Y = 51 else
"111111111111" when X = 224 AND Y = 51 else
"111111111111" when X = 225 AND Y = 51 else
"111111111111" when X = 226 AND Y = 51 else
"111111111111" when X = 227 AND Y = 51 else
"111111111111" when X = 228 AND Y = 51 else
"111111111111" when X = 229 AND Y = 51 else
"111111111111" when X = 230 AND Y = 51 else
"111111111111" when X = 231 AND Y = 51 else
"111111111111" when X = 232 AND Y = 51 else
"111111111111" when X = 233 AND Y = 51 else
"111111111111" when X = 234 AND Y = 51 else
"111111111111" when X = 235 AND Y = 51 else
"111111111111" when X = 236 AND Y = 51 else
"111111111111" when X = 237 AND Y = 51 else
"111111111111" when X = 238 AND Y = 51 else
"111111111111" when X = 239 AND Y = 51 else
"111111111111" when X = 240 AND Y = 51 else
"111111111111" when X = 241 AND Y = 51 else
"111111111111" when X = 242 AND Y = 51 else
"111111111111" when X = 243 AND Y = 51 else
"111111111111" when X = 244 AND Y = 51 else
"111111111111" when X = 245 AND Y = 51 else
"111111111111" when X = 246 AND Y = 51 else
"111111111111" when X = 247 AND Y = 51 else
"111111111111" when X = 248 AND Y = 51 else
"111111111111" when X = 249 AND Y = 51 else
"111111111111" when X = 250 AND Y = 51 else
"111111111111" when X = 251 AND Y = 51 else
"111111111111" when X = 252 AND Y = 51 else
"111111111111" when X = 253 AND Y = 51 else
"111111111111" when X = 254 AND Y = 51 else
"111111111111" when X = 255 AND Y = 51 else
"111111111111" when X = 256 AND Y = 51 else
"111111111111" when X = 257 AND Y = 51 else
"111111111111" when X = 258 AND Y = 51 else
"111111111111" when X = 259 AND Y = 51 else
"111111111111" when X = 260 AND Y = 51 else
"111111111111" when X = 261 AND Y = 51 else
"111111111111" when X = 262 AND Y = 51 else
"111111111111" when X = 263 AND Y = 51 else
"111111111111" when X = 264 AND Y = 51 else
"110111011111" when X = 265 AND Y = 51 else
"110111011111" when X = 266 AND Y = 51 else
"110111011111" when X = 267 AND Y = 51 else
"110111011111" when X = 268 AND Y = 51 else
"110111011111" when X = 269 AND Y = 51 else
"110111011111" when X = 270 AND Y = 51 else
"110111011111" when X = 271 AND Y = 51 else
"110111011111" when X = 272 AND Y = 51 else
"110111011111" when X = 273 AND Y = 51 else
"110111011111" when X = 274 AND Y = 51 else
"110111011111" when X = 275 AND Y = 51 else
"110111011111" when X = 276 AND Y = 51 else
"110111011111" when X = 277 AND Y = 51 else
"110111011111" when X = 278 AND Y = 51 else
"110111011111" when X = 279 AND Y = 51 else
"000000000000" when X = 280 AND Y = 51 else
"000000000000" when X = 281 AND Y = 51 else
"000000000000" when X = 282 AND Y = 51 else
"000000000000" when X = 283 AND Y = 51 else
"000000000000" when X = 284 AND Y = 51 else
"000000000000" when X = 285 AND Y = 51 else
"000000000000" when X = 286 AND Y = 51 else
"000000000000" when X = 287 AND Y = 51 else
"000000000000" when X = 288 AND Y = 51 else
"000000000000" when X = 289 AND Y = 51 else
"000000000000" when X = 290 AND Y = 51 else
"000000000000" when X = 291 AND Y = 51 else
"000000000000" when X = 292 AND Y = 51 else
"000000000000" when X = 293 AND Y = 51 else
"000000000000" when X = 294 AND Y = 51 else
"000000000000" when X = 295 AND Y = 51 else
"000000000000" when X = 296 AND Y = 51 else
"000000000000" when X = 297 AND Y = 51 else
"000000000000" when X = 298 AND Y = 51 else
"000000000000" when X = 299 AND Y = 51 else
"000000000000" when X = 300 AND Y = 51 else
"000000000000" when X = 301 AND Y = 51 else
"000000000000" when X = 302 AND Y = 51 else
"000000000000" when X = 303 AND Y = 51 else
"000000000000" when X = 304 AND Y = 51 else
"000000000000" when X = 305 AND Y = 51 else
"000000000000" when X = 306 AND Y = 51 else
"000000000000" when X = 307 AND Y = 51 else
"000000000000" when X = 308 AND Y = 51 else
"000000000000" when X = 309 AND Y = 51 else
"000000000000" when X = 310 AND Y = 51 else
"000000000000" when X = 311 AND Y = 51 else
"000000000000" when X = 312 AND Y = 51 else
"000000000000" when X = 313 AND Y = 51 else
"000000000000" when X = 314 AND Y = 51 else
"000000000000" when X = 315 AND Y = 51 else
"000000000000" when X = 316 AND Y = 51 else
"000000000000" when X = 317 AND Y = 51 else
"000000000000" when X = 318 AND Y = 51 else
"000000000000" when X = 319 AND Y = 51 else
"000000000000" when X = 320 AND Y = 51 else
"000000000000" when X = 321 AND Y = 51 else
"000000000000" when X = 322 AND Y = 51 else
"000000000000" when X = 323 AND Y = 51 else
"000000000000" when X = 324 AND Y = 51 else
"100010011101" when X = 0 AND Y = 52 else
"100010011101" when X = 1 AND Y = 52 else
"100010011101" when X = 2 AND Y = 52 else
"100010011101" when X = 3 AND Y = 52 else
"100010011101" when X = 4 AND Y = 52 else
"100010011101" when X = 5 AND Y = 52 else
"100010011101" when X = 6 AND Y = 52 else
"100010011101" when X = 7 AND Y = 52 else
"100010011101" when X = 8 AND Y = 52 else
"100010011101" when X = 9 AND Y = 52 else
"100010011101" when X = 10 AND Y = 52 else
"100010011101" when X = 11 AND Y = 52 else
"100010011101" when X = 12 AND Y = 52 else
"100010011101" when X = 13 AND Y = 52 else
"100010011101" when X = 14 AND Y = 52 else
"100010011101" when X = 15 AND Y = 52 else
"100010011101" when X = 16 AND Y = 52 else
"100010011101" when X = 17 AND Y = 52 else
"100010011101" when X = 18 AND Y = 52 else
"100010011101" when X = 19 AND Y = 52 else
"100010011101" when X = 20 AND Y = 52 else
"100010011101" when X = 21 AND Y = 52 else
"100010011101" when X = 22 AND Y = 52 else
"100010011101" when X = 23 AND Y = 52 else
"100010011101" when X = 24 AND Y = 52 else
"100010011101" when X = 25 AND Y = 52 else
"100010011101" when X = 26 AND Y = 52 else
"100010011101" when X = 27 AND Y = 52 else
"100010011101" when X = 28 AND Y = 52 else
"100010011101" when X = 29 AND Y = 52 else
"100010011101" when X = 30 AND Y = 52 else
"100010011101" when X = 31 AND Y = 52 else
"100010011101" when X = 32 AND Y = 52 else
"100010011101" when X = 33 AND Y = 52 else
"100010011101" when X = 34 AND Y = 52 else
"100010011101" when X = 35 AND Y = 52 else
"100010011101" when X = 36 AND Y = 52 else
"100010011101" when X = 37 AND Y = 52 else
"100010011101" when X = 38 AND Y = 52 else
"100010011101" when X = 39 AND Y = 52 else
"100010011101" when X = 40 AND Y = 52 else
"100010011101" when X = 41 AND Y = 52 else
"100010011101" when X = 42 AND Y = 52 else
"100010011101" when X = 43 AND Y = 52 else
"100010011101" when X = 44 AND Y = 52 else
"110111011111" when X = 45 AND Y = 52 else
"110111011111" when X = 46 AND Y = 52 else
"110111011111" when X = 47 AND Y = 52 else
"110111011111" when X = 48 AND Y = 52 else
"110111011111" when X = 49 AND Y = 52 else
"110111011111" when X = 50 AND Y = 52 else
"110111011111" when X = 51 AND Y = 52 else
"110111011111" when X = 52 AND Y = 52 else
"110111011111" when X = 53 AND Y = 52 else
"110111011111" when X = 54 AND Y = 52 else
"110111011111" when X = 55 AND Y = 52 else
"110111011111" when X = 56 AND Y = 52 else
"110111011111" when X = 57 AND Y = 52 else
"110111011111" when X = 58 AND Y = 52 else
"110111011111" when X = 59 AND Y = 52 else
"110111011111" when X = 60 AND Y = 52 else
"110111011111" when X = 61 AND Y = 52 else
"110111011111" when X = 62 AND Y = 52 else
"110111011111" when X = 63 AND Y = 52 else
"110111011111" when X = 64 AND Y = 52 else
"110111011111" when X = 65 AND Y = 52 else
"110111011111" when X = 66 AND Y = 52 else
"110111011111" when X = 67 AND Y = 52 else
"110111011111" when X = 68 AND Y = 52 else
"110111011111" when X = 69 AND Y = 52 else
"111111111111" when X = 70 AND Y = 52 else
"111111111111" when X = 71 AND Y = 52 else
"111111111111" when X = 72 AND Y = 52 else
"111111111111" when X = 73 AND Y = 52 else
"111111111111" when X = 74 AND Y = 52 else
"111111111111" when X = 75 AND Y = 52 else
"111111111111" when X = 76 AND Y = 52 else
"111111111111" when X = 77 AND Y = 52 else
"111111111111" when X = 78 AND Y = 52 else
"111111111111" when X = 79 AND Y = 52 else
"111111111111" when X = 80 AND Y = 52 else
"111111111111" when X = 81 AND Y = 52 else
"111111111111" when X = 82 AND Y = 52 else
"111111111111" when X = 83 AND Y = 52 else
"111111111111" when X = 84 AND Y = 52 else
"111111111111" when X = 85 AND Y = 52 else
"111111111111" when X = 86 AND Y = 52 else
"111111111111" when X = 87 AND Y = 52 else
"111111111111" when X = 88 AND Y = 52 else
"111111111111" when X = 89 AND Y = 52 else
"111111111111" when X = 90 AND Y = 52 else
"111111111111" when X = 91 AND Y = 52 else
"111111111111" when X = 92 AND Y = 52 else
"111111111111" when X = 93 AND Y = 52 else
"111111111111" when X = 94 AND Y = 52 else
"111111111111" when X = 95 AND Y = 52 else
"111111111111" when X = 96 AND Y = 52 else
"111111111111" when X = 97 AND Y = 52 else
"111111111111" when X = 98 AND Y = 52 else
"111111111111" when X = 99 AND Y = 52 else
"111111111111" when X = 100 AND Y = 52 else
"111111111111" when X = 101 AND Y = 52 else
"111111111111" when X = 102 AND Y = 52 else
"111111111111" when X = 103 AND Y = 52 else
"111111111111" when X = 104 AND Y = 52 else
"111111111111" when X = 105 AND Y = 52 else
"111111111111" when X = 106 AND Y = 52 else
"111111111111" when X = 107 AND Y = 52 else
"111111111111" when X = 108 AND Y = 52 else
"111111111111" when X = 109 AND Y = 52 else
"111111111111" when X = 110 AND Y = 52 else
"111111111111" when X = 111 AND Y = 52 else
"111111111111" when X = 112 AND Y = 52 else
"111111111111" when X = 113 AND Y = 52 else
"111111111111" when X = 114 AND Y = 52 else
"111111111111" when X = 115 AND Y = 52 else
"111111111111" when X = 116 AND Y = 52 else
"111111111111" when X = 117 AND Y = 52 else
"111111111111" when X = 118 AND Y = 52 else
"111111111111" when X = 119 AND Y = 52 else
"111111111111" when X = 120 AND Y = 52 else
"111111111111" when X = 121 AND Y = 52 else
"111111111111" when X = 122 AND Y = 52 else
"111111111111" when X = 123 AND Y = 52 else
"111111111111" when X = 124 AND Y = 52 else
"111111111111" when X = 125 AND Y = 52 else
"111111111111" when X = 126 AND Y = 52 else
"111111111111" when X = 127 AND Y = 52 else
"111111111111" when X = 128 AND Y = 52 else
"111111111111" when X = 129 AND Y = 52 else
"111111111111" when X = 130 AND Y = 52 else
"111111111111" when X = 131 AND Y = 52 else
"111111111111" when X = 132 AND Y = 52 else
"111111111111" when X = 133 AND Y = 52 else
"111111111111" when X = 134 AND Y = 52 else
"111111111111" when X = 135 AND Y = 52 else
"111111111111" when X = 136 AND Y = 52 else
"111111111111" when X = 137 AND Y = 52 else
"111111111111" when X = 138 AND Y = 52 else
"111111111111" when X = 139 AND Y = 52 else
"111111111111" when X = 140 AND Y = 52 else
"111111111111" when X = 141 AND Y = 52 else
"111111111111" when X = 142 AND Y = 52 else
"111111111111" when X = 143 AND Y = 52 else
"111111111111" when X = 144 AND Y = 52 else
"111111111111" when X = 145 AND Y = 52 else
"111111111111" when X = 146 AND Y = 52 else
"111111111111" when X = 147 AND Y = 52 else
"111111111111" when X = 148 AND Y = 52 else
"111111111111" when X = 149 AND Y = 52 else
"111111111111" when X = 150 AND Y = 52 else
"111111111111" when X = 151 AND Y = 52 else
"111111111111" when X = 152 AND Y = 52 else
"111111111111" when X = 153 AND Y = 52 else
"111111111111" when X = 154 AND Y = 52 else
"111111111111" when X = 155 AND Y = 52 else
"111111111111" when X = 156 AND Y = 52 else
"111111111111" when X = 157 AND Y = 52 else
"111111111111" when X = 158 AND Y = 52 else
"111111111111" when X = 159 AND Y = 52 else
"111111111111" when X = 160 AND Y = 52 else
"111111111111" when X = 161 AND Y = 52 else
"111111111111" when X = 162 AND Y = 52 else
"111111111111" when X = 163 AND Y = 52 else
"111111111111" when X = 164 AND Y = 52 else
"111111111111" when X = 165 AND Y = 52 else
"111111111111" when X = 166 AND Y = 52 else
"111111111111" when X = 167 AND Y = 52 else
"111111111111" when X = 168 AND Y = 52 else
"111111111111" when X = 169 AND Y = 52 else
"111111111111" when X = 170 AND Y = 52 else
"111111111111" when X = 171 AND Y = 52 else
"111111111111" when X = 172 AND Y = 52 else
"111111111111" when X = 173 AND Y = 52 else
"111111111111" when X = 174 AND Y = 52 else
"111111111111" when X = 175 AND Y = 52 else
"111111111111" when X = 176 AND Y = 52 else
"111111111111" when X = 177 AND Y = 52 else
"111111111111" when X = 178 AND Y = 52 else
"111111111111" when X = 179 AND Y = 52 else
"111111111111" when X = 180 AND Y = 52 else
"111111111111" when X = 181 AND Y = 52 else
"111111111111" when X = 182 AND Y = 52 else
"111111111111" when X = 183 AND Y = 52 else
"111111111111" when X = 184 AND Y = 52 else
"111111111111" when X = 185 AND Y = 52 else
"111111111111" when X = 186 AND Y = 52 else
"111111111111" when X = 187 AND Y = 52 else
"111111111111" when X = 188 AND Y = 52 else
"111111111111" when X = 189 AND Y = 52 else
"111111111111" when X = 190 AND Y = 52 else
"111111111111" when X = 191 AND Y = 52 else
"111111111111" when X = 192 AND Y = 52 else
"111111111111" when X = 193 AND Y = 52 else
"111111111111" when X = 194 AND Y = 52 else
"111111111111" when X = 195 AND Y = 52 else
"111111111111" when X = 196 AND Y = 52 else
"111111111111" when X = 197 AND Y = 52 else
"111111111111" when X = 198 AND Y = 52 else
"111111111111" when X = 199 AND Y = 52 else
"111111111111" when X = 200 AND Y = 52 else
"111111111111" when X = 201 AND Y = 52 else
"111111111111" when X = 202 AND Y = 52 else
"111111111111" when X = 203 AND Y = 52 else
"111111111111" when X = 204 AND Y = 52 else
"111111111111" when X = 205 AND Y = 52 else
"111111111111" when X = 206 AND Y = 52 else
"111111111111" when X = 207 AND Y = 52 else
"111111111111" when X = 208 AND Y = 52 else
"111111111111" when X = 209 AND Y = 52 else
"111111111111" when X = 210 AND Y = 52 else
"111111111111" when X = 211 AND Y = 52 else
"111111111111" when X = 212 AND Y = 52 else
"111111111111" when X = 213 AND Y = 52 else
"111111111111" when X = 214 AND Y = 52 else
"111111111111" when X = 215 AND Y = 52 else
"111111111111" when X = 216 AND Y = 52 else
"111111111111" when X = 217 AND Y = 52 else
"111111111111" when X = 218 AND Y = 52 else
"111111111111" when X = 219 AND Y = 52 else
"111111111111" when X = 220 AND Y = 52 else
"111111111111" when X = 221 AND Y = 52 else
"111111111111" when X = 222 AND Y = 52 else
"111111111111" when X = 223 AND Y = 52 else
"111111111111" when X = 224 AND Y = 52 else
"111111111111" when X = 225 AND Y = 52 else
"111111111111" when X = 226 AND Y = 52 else
"111111111111" when X = 227 AND Y = 52 else
"111111111111" when X = 228 AND Y = 52 else
"111111111111" when X = 229 AND Y = 52 else
"111111111111" when X = 230 AND Y = 52 else
"111111111111" when X = 231 AND Y = 52 else
"111111111111" when X = 232 AND Y = 52 else
"111111111111" when X = 233 AND Y = 52 else
"111111111111" when X = 234 AND Y = 52 else
"111111111111" when X = 235 AND Y = 52 else
"111111111111" when X = 236 AND Y = 52 else
"111111111111" when X = 237 AND Y = 52 else
"111111111111" when X = 238 AND Y = 52 else
"111111111111" when X = 239 AND Y = 52 else
"111111111111" when X = 240 AND Y = 52 else
"111111111111" when X = 241 AND Y = 52 else
"111111111111" when X = 242 AND Y = 52 else
"111111111111" when X = 243 AND Y = 52 else
"111111111111" when X = 244 AND Y = 52 else
"111111111111" when X = 245 AND Y = 52 else
"111111111111" when X = 246 AND Y = 52 else
"111111111111" when X = 247 AND Y = 52 else
"111111111111" when X = 248 AND Y = 52 else
"111111111111" when X = 249 AND Y = 52 else
"111111111111" when X = 250 AND Y = 52 else
"111111111111" when X = 251 AND Y = 52 else
"111111111111" when X = 252 AND Y = 52 else
"111111111111" when X = 253 AND Y = 52 else
"111111111111" when X = 254 AND Y = 52 else
"111111111111" when X = 255 AND Y = 52 else
"111111111111" when X = 256 AND Y = 52 else
"111111111111" when X = 257 AND Y = 52 else
"111111111111" when X = 258 AND Y = 52 else
"111111111111" when X = 259 AND Y = 52 else
"111111111111" when X = 260 AND Y = 52 else
"111111111111" when X = 261 AND Y = 52 else
"111111111111" when X = 262 AND Y = 52 else
"111111111111" when X = 263 AND Y = 52 else
"111111111111" when X = 264 AND Y = 52 else
"110111011111" when X = 265 AND Y = 52 else
"110111011111" when X = 266 AND Y = 52 else
"110111011111" when X = 267 AND Y = 52 else
"110111011111" when X = 268 AND Y = 52 else
"110111011111" when X = 269 AND Y = 52 else
"110111011111" when X = 270 AND Y = 52 else
"110111011111" when X = 271 AND Y = 52 else
"110111011111" when X = 272 AND Y = 52 else
"110111011111" when X = 273 AND Y = 52 else
"110111011111" when X = 274 AND Y = 52 else
"110111011111" when X = 275 AND Y = 52 else
"110111011111" when X = 276 AND Y = 52 else
"110111011111" when X = 277 AND Y = 52 else
"110111011111" when X = 278 AND Y = 52 else
"110111011111" when X = 279 AND Y = 52 else
"000000000000" when X = 280 AND Y = 52 else
"000000000000" when X = 281 AND Y = 52 else
"000000000000" when X = 282 AND Y = 52 else
"000000000000" when X = 283 AND Y = 52 else
"000000000000" when X = 284 AND Y = 52 else
"000000000000" when X = 285 AND Y = 52 else
"000000000000" when X = 286 AND Y = 52 else
"000000000000" when X = 287 AND Y = 52 else
"000000000000" when X = 288 AND Y = 52 else
"000000000000" when X = 289 AND Y = 52 else
"000000000000" when X = 290 AND Y = 52 else
"000000000000" when X = 291 AND Y = 52 else
"000000000000" when X = 292 AND Y = 52 else
"000000000000" when X = 293 AND Y = 52 else
"000000000000" when X = 294 AND Y = 52 else
"000000000000" when X = 295 AND Y = 52 else
"000000000000" when X = 296 AND Y = 52 else
"000000000000" when X = 297 AND Y = 52 else
"000000000000" when X = 298 AND Y = 52 else
"000000000000" when X = 299 AND Y = 52 else
"000000000000" when X = 300 AND Y = 52 else
"000000000000" when X = 301 AND Y = 52 else
"000000000000" when X = 302 AND Y = 52 else
"000000000000" when X = 303 AND Y = 52 else
"000000000000" when X = 304 AND Y = 52 else
"000000000000" when X = 305 AND Y = 52 else
"000000000000" when X = 306 AND Y = 52 else
"000000000000" when X = 307 AND Y = 52 else
"000000000000" when X = 308 AND Y = 52 else
"000000000000" when X = 309 AND Y = 52 else
"000000000000" when X = 310 AND Y = 52 else
"000000000000" when X = 311 AND Y = 52 else
"000000000000" when X = 312 AND Y = 52 else
"000000000000" when X = 313 AND Y = 52 else
"000000000000" when X = 314 AND Y = 52 else
"000000000000" when X = 315 AND Y = 52 else
"000000000000" when X = 316 AND Y = 52 else
"000000000000" when X = 317 AND Y = 52 else
"000000000000" when X = 318 AND Y = 52 else
"000000000000" when X = 319 AND Y = 52 else
"000000000000" when X = 320 AND Y = 52 else
"000000000000" when X = 321 AND Y = 52 else
"000000000000" when X = 322 AND Y = 52 else
"000000000000" when X = 323 AND Y = 52 else
"000000000000" when X = 324 AND Y = 52 else
"100010011101" when X = 0 AND Y = 53 else
"100010011101" when X = 1 AND Y = 53 else
"100010011101" when X = 2 AND Y = 53 else
"100010011101" when X = 3 AND Y = 53 else
"100010011101" when X = 4 AND Y = 53 else
"100010011101" when X = 5 AND Y = 53 else
"100010011101" when X = 6 AND Y = 53 else
"100010011101" when X = 7 AND Y = 53 else
"100010011101" when X = 8 AND Y = 53 else
"100010011101" when X = 9 AND Y = 53 else
"100010011101" when X = 10 AND Y = 53 else
"100010011101" when X = 11 AND Y = 53 else
"100010011101" when X = 12 AND Y = 53 else
"100010011101" when X = 13 AND Y = 53 else
"100010011101" when X = 14 AND Y = 53 else
"100010011101" when X = 15 AND Y = 53 else
"100010011101" when X = 16 AND Y = 53 else
"100010011101" when X = 17 AND Y = 53 else
"100010011101" when X = 18 AND Y = 53 else
"100010011101" when X = 19 AND Y = 53 else
"100010011101" when X = 20 AND Y = 53 else
"100010011101" when X = 21 AND Y = 53 else
"100010011101" when X = 22 AND Y = 53 else
"100010011101" when X = 23 AND Y = 53 else
"100010011101" when X = 24 AND Y = 53 else
"100010011101" when X = 25 AND Y = 53 else
"100010011101" when X = 26 AND Y = 53 else
"100010011101" when X = 27 AND Y = 53 else
"100010011101" when X = 28 AND Y = 53 else
"100010011101" when X = 29 AND Y = 53 else
"100010011101" when X = 30 AND Y = 53 else
"100010011101" when X = 31 AND Y = 53 else
"100010011101" when X = 32 AND Y = 53 else
"100010011101" when X = 33 AND Y = 53 else
"100010011101" when X = 34 AND Y = 53 else
"100010011101" when X = 35 AND Y = 53 else
"100010011101" when X = 36 AND Y = 53 else
"100010011101" when X = 37 AND Y = 53 else
"100010011101" when X = 38 AND Y = 53 else
"100010011101" when X = 39 AND Y = 53 else
"100010011101" when X = 40 AND Y = 53 else
"100010011101" when X = 41 AND Y = 53 else
"100010011101" when X = 42 AND Y = 53 else
"100010011101" when X = 43 AND Y = 53 else
"100010011101" when X = 44 AND Y = 53 else
"110111011111" when X = 45 AND Y = 53 else
"110111011111" when X = 46 AND Y = 53 else
"110111011111" when X = 47 AND Y = 53 else
"110111011111" when X = 48 AND Y = 53 else
"110111011111" when X = 49 AND Y = 53 else
"110111011111" when X = 50 AND Y = 53 else
"110111011111" when X = 51 AND Y = 53 else
"110111011111" when X = 52 AND Y = 53 else
"110111011111" when X = 53 AND Y = 53 else
"110111011111" when X = 54 AND Y = 53 else
"110111011111" when X = 55 AND Y = 53 else
"110111011111" when X = 56 AND Y = 53 else
"110111011111" when X = 57 AND Y = 53 else
"110111011111" when X = 58 AND Y = 53 else
"110111011111" when X = 59 AND Y = 53 else
"110111011111" when X = 60 AND Y = 53 else
"110111011111" when X = 61 AND Y = 53 else
"110111011111" when X = 62 AND Y = 53 else
"110111011111" when X = 63 AND Y = 53 else
"110111011111" when X = 64 AND Y = 53 else
"110111011111" when X = 65 AND Y = 53 else
"110111011111" when X = 66 AND Y = 53 else
"110111011111" when X = 67 AND Y = 53 else
"110111011111" when X = 68 AND Y = 53 else
"110111011111" when X = 69 AND Y = 53 else
"111111111111" when X = 70 AND Y = 53 else
"111111111111" when X = 71 AND Y = 53 else
"111111111111" when X = 72 AND Y = 53 else
"111111111111" when X = 73 AND Y = 53 else
"111111111111" when X = 74 AND Y = 53 else
"111111111111" when X = 75 AND Y = 53 else
"111111111111" when X = 76 AND Y = 53 else
"111111111111" when X = 77 AND Y = 53 else
"111111111111" when X = 78 AND Y = 53 else
"111111111111" when X = 79 AND Y = 53 else
"111111111111" when X = 80 AND Y = 53 else
"111111111111" when X = 81 AND Y = 53 else
"111111111111" when X = 82 AND Y = 53 else
"111111111111" when X = 83 AND Y = 53 else
"111111111111" when X = 84 AND Y = 53 else
"111111111111" when X = 85 AND Y = 53 else
"111111111111" when X = 86 AND Y = 53 else
"111111111111" when X = 87 AND Y = 53 else
"111111111111" when X = 88 AND Y = 53 else
"111111111111" when X = 89 AND Y = 53 else
"111111111111" when X = 90 AND Y = 53 else
"111111111111" when X = 91 AND Y = 53 else
"111111111111" when X = 92 AND Y = 53 else
"111111111111" when X = 93 AND Y = 53 else
"111111111111" when X = 94 AND Y = 53 else
"111111111111" when X = 95 AND Y = 53 else
"111111111111" when X = 96 AND Y = 53 else
"111111111111" when X = 97 AND Y = 53 else
"111111111111" when X = 98 AND Y = 53 else
"111111111111" when X = 99 AND Y = 53 else
"111111111111" when X = 100 AND Y = 53 else
"111111111111" when X = 101 AND Y = 53 else
"111111111111" when X = 102 AND Y = 53 else
"111111111111" when X = 103 AND Y = 53 else
"111111111111" when X = 104 AND Y = 53 else
"111111111111" when X = 105 AND Y = 53 else
"111111111111" when X = 106 AND Y = 53 else
"111111111111" when X = 107 AND Y = 53 else
"111111111111" when X = 108 AND Y = 53 else
"111111111111" when X = 109 AND Y = 53 else
"111111111111" when X = 110 AND Y = 53 else
"111111111111" when X = 111 AND Y = 53 else
"111111111111" when X = 112 AND Y = 53 else
"111111111111" when X = 113 AND Y = 53 else
"111111111111" when X = 114 AND Y = 53 else
"111111111111" when X = 115 AND Y = 53 else
"111111111111" when X = 116 AND Y = 53 else
"111111111111" when X = 117 AND Y = 53 else
"111111111111" when X = 118 AND Y = 53 else
"111111111111" when X = 119 AND Y = 53 else
"111111111111" when X = 120 AND Y = 53 else
"111111111111" when X = 121 AND Y = 53 else
"111111111111" when X = 122 AND Y = 53 else
"111111111111" when X = 123 AND Y = 53 else
"111111111111" when X = 124 AND Y = 53 else
"111111111111" when X = 125 AND Y = 53 else
"111111111111" when X = 126 AND Y = 53 else
"111111111111" when X = 127 AND Y = 53 else
"111111111111" when X = 128 AND Y = 53 else
"111111111111" when X = 129 AND Y = 53 else
"111111111111" when X = 130 AND Y = 53 else
"111111111111" when X = 131 AND Y = 53 else
"111111111111" when X = 132 AND Y = 53 else
"111111111111" when X = 133 AND Y = 53 else
"111111111111" when X = 134 AND Y = 53 else
"111111111111" when X = 135 AND Y = 53 else
"111111111111" when X = 136 AND Y = 53 else
"111111111111" when X = 137 AND Y = 53 else
"111111111111" when X = 138 AND Y = 53 else
"111111111111" when X = 139 AND Y = 53 else
"111111111111" when X = 140 AND Y = 53 else
"111111111111" when X = 141 AND Y = 53 else
"111111111111" when X = 142 AND Y = 53 else
"111111111111" when X = 143 AND Y = 53 else
"111111111111" when X = 144 AND Y = 53 else
"111111111111" when X = 145 AND Y = 53 else
"111111111111" when X = 146 AND Y = 53 else
"111111111111" when X = 147 AND Y = 53 else
"111111111111" when X = 148 AND Y = 53 else
"111111111111" when X = 149 AND Y = 53 else
"111111111111" when X = 150 AND Y = 53 else
"111111111111" when X = 151 AND Y = 53 else
"111111111111" when X = 152 AND Y = 53 else
"111111111111" when X = 153 AND Y = 53 else
"111111111111" when X = 154 AND Y = 53 else
"111111111111" when X = 155 AND Y = 53 else
"111111111111" when X = 156 AND Y = 53 else
"111111111111" when X = 157 AND Y = 53 else
"111111111111" when X = 158 AND Y = 53 else
"111111111111" when X = 159 AND Y = 53 else
"111111111111" when X = 160 AND Y = 53 else
"111111111111" when X = 161 AND Y = 53 else
"111111111111" when X = 162 AND Y = 53 else
"111111111111" when X = 163 AND Y = 53 else
"111111111111" when X = 164 AND Y = 53 else
"111111111111" when X = 165 AND Y = 53 else
"111111111111" when X = 166 AND Y = 53 else
"111111111111" when X = 167 AND Y = 53 else
"111111111111" when X = 168 AND Y = 53 else
"111111111111" when X = 169 AND Y = 53 else
"111111111111" when X = 170 AND Y = 53 else
"111111111111" when X = 171 AND Y = 53 else
"111111111111" when X = 172 AND Y = 53 else
"111111111111" when X = 173 AND Y = 53 else
"111111111111" when X = 174 AND Y = 53 else
"111111111111" when X = 175 AND Y = 53 else
"111111111111" when X = 176 AND Y = 53 else
"111111111111" when X = 177 AND Y = 53 else
"111111111111" when X = 178 AND Y = 53 else
"111111111111" when X = 179 AND Y = 53 else
"111111111111" when X = 180 AND Y = 53 else
"111111111111" when X = 181 AND Y = 53 else
"111111111111" when X = 182 AND Y = 53 else
"111111111111" when X = 183 AND Y = 53 else
"111111111111" when X = 184 AND Y = 53 else
"111111111111" when X = 185 AND Y = 53 else
"111111111111" when X = 186 AND Y = 53 else
"111111111111" when X = 187 AND Y = 53 else
"111111111111" when X = 188 AND Y = 53 else
"111111111111" when X = 189 AND Y = 53 else
"111111111111" when X = 190 AND Y = 53 else
"111111111111" when X = 191 AND Y = 53 else
"111111111111" when X = 192 AND Y = 53 else
"111111111111" when X = 193 AND Y = 53 else
"111111111111" when X = 194 AND Y = 53 else
"111111111111" when X = 195 AND Y = 53 else
"111111111111" when X = 196 AND Y = 53 else
"111111111111" when X = 197 AND Y = 53 else
"111111111111" when X = 198 AND Y = 53 else
"111111111111" when X = 199 AND Y = 53 else
"111111111111" when X = 200 AND Y = 53 else
"111111111111" when X = 201 AND Y = 53 else
"111111111111" when X = 202 AND Y = 53 else
"111111111111" when X = 203 AND Y = 53 else
"111111111111" when X = 204 AND Y = 53 else
"111111111111" when X = 205 AND Y = 53 else
"111111111111" when X = 206 AND Y = 53 else
"111111111111" when X = 207 AND Y = 53 else
"111111111111" when X = 208 AND Y = 53 else
"111111111111" when X = 209 AND Y = 53 else
"111111111111" when X = 210 AND Y = 53 else
"111111111111" when X = 211 AND Y = 53 else
"111111111111" when X = 212 AND Y = 53 else
"111111111111" when X = 213 AND Y = 53 else
"111111111111" when X = 214 AND Y = 53 else
"111111111111" when X = 215 AND Y = 53 else
"111111111111" when X = 216 AND Y = 53 else
"111111111111" when X = 217 AND Y = 53 else
"111111111111" when X = 218 AND Y = 53 else
"111111111111" when X = 219 AND Y = 53 else
"111111111111" when X = 220 AND Y = 53 else
"111111111111" when X = 221 AND Y = 53 else
"111111111111" when X = 222 AND Y = 53 else
"111111111111" when X = 223 AND Y = 53 else
"111111111111" when X = 224 AND Y = 53 else
"111111111111" when X = 225 AND Y = 53 else
"111111111111" when X = 226 AND Y = 53 else
"111111111111" when X = 227 AND Y = 53 else
"111111111111" when X = 228 AND Y = 53 else
"111111111111" when X = 229 AND Y = 53 else
"111111111111" when X = 230 AND Y = 53 else
"111111111111" when X = 231 AND Y = 53 else
"111111111111" when X = 232 AND Y = 53 else
"111111111111" when X = 233 AND Y = 53 else
"111111111111" when X = 234 AND Y = 53 else
"111111111111" when X = 235 AND Y = 53 else
"111111111111" when X = 236 AND Y = 53 else
"111111111111" when X = 237 AND Y = 53 else
"111111111111" when X = 238 AND Y = 53 else
"111111111111" when X = 239 AND Y = 53 else
"111111111111" when X = 240 AND Y = 53 else
"111111111111" when X = 241 AND Y = 53 else
"111111111111" when X = 242 AND Y = 53 else
"111111111111" when X = 243 AND Y = 53 else
"111111111111" when X = 244 AND Y = 53 else
"111111111111" when X = 245 AND Y = 53 else
"111111111111" when X = 246 AND Y = 53 else
"111111111111" when X = 247 AND Y = 53 else
"111111111111" when X = 248 AND Y = 53 else
"111111111111" when X = 249 AND Y = 53 else
"111111111111" when X = 250 AND Y = 53 else
"111111111111" when X = 251 AND Y = 53 else
"111111111111" when X = 252 AND Y = 53 else
"111111111111" when X = 253 AND Y = 53 else
"111111111111" when X = 254 AND Y = 53 else
"111111111111" when X = 255 AND Y = 53 else
"111111111111" when X = 256 AND Y = 53 else
"111111111111" when X = 257 AND Y = 53 else
"111111111111" when X = 258 AND Y = 53 else
"111111111111" when X = 259 AND Y = 53 else
"111111111111" when X = 260 AND Y = 53 else
"111111111111" when X = 261 AND Y = 53 else
"111111111111" when X = 262 AND Y = 53 else
"111111111111" when X = 263 AND Y = 53 else
"111111111111" when X = 264 AND Y = 53 else
"110111011111" when X = 265 AND Y = 53 else
"110111011111" when X = 266 AND Y = 53 else
"110111011111" when X = 267 AND Y = 53 else
"110111011111" when X = 268 AND Y = 53 else
"110111011111" when X = 269 AND Y = 53 else
"110111011111" when X = 270 AND Y = 53 else
"110111011111" when X = 271 AND Y = 53 else
"110111011111" when X = 272 AND Y = 53 else
"110111011111" when X = 273 AND Y = 53 else
"110111011111" when X = 274 AND Y = 53 else
"110111011111" when X = 275 AND Y = 53 else
"110111011111" when X = 276 AND Y = 53 else
"110111011111" when X = 277 AND Y = 53 else
"110111011111" when X = 278 AND Y = 53 else
"110111011111" when X = 279 AND Y = 53 else
"000000000000" when X = 280 AND Y = 53 else
"000000000000" when X = 281 AND Y = 53 else
"000000000000" when X = 282 AND Y = 53 else
"000000000000" when X = 283 AND Y = 53 else
"000000000000" when X = 284 AND Y = 53 else
"000000000000" when X = 285 AND Y = 53 else
"000000000000" when X = 286 AND Y = 53 else
"000000000000" when X = 287 AND Y = 53 else
"000000000000" when X = 288 AND Y = 53 else
"000000000000" when X = 289 AND Y = 53 else
"000000000000" when X = 290 AND Y = 53 else
"000000000000" when X = 291 AND Y = 53 else
"000000000000" when X = 292 AND Y = 53 else
"000000000000" when X = 293 AND Y = 53 else
"000000000000" when X = 294 AND Y = 53 else
"000000000000" when X = 295 AND Y = 53 else
"000000000000" when X = 296 AND Y = 53 else
"000000000000" when X = 297 AND Y = 53 else
"000000000000" when X = 298 AND Y = 53 else
"000000000000" when X = 299 AND Y = 53 else
"000000000000" when X = 300 AND Y = 53 else
"000000000000" when X = 301 AND Y = 53 else
"000000000000" when X = 302 AND Y = 53 else
"000000000000" when X = 303 AND Y = 53 else
"000000000000" when X = 304 AND Y = 53 else
"000000000000" when X = 305 AND Y = 53 else
"000000000000" when X = 306 AND Y = 53 else
"000000000000" when X = 307 AND Y = 53 else
"000000000000" when X = 308 AND Y = 53 else
"000000000000" when X = 309 AND Y = 53 else
"000000000000" when X = 310 AND Y = 53 else
"000000000000" when X = 311 AND Y = 53 else
"000000000000" when X = 312 AND Y = 53 else
"000000000000" when X = 313 AND Y = 53 else
"000000000000" when X = 314 AND Y = 53 else
"000000000000" when X = 315 AND Y = 53 else
"000000000000" when X = 316 AND Y = 53 else
"000000000000" when X = 317 AND Y = 53 else
"000000000000" when X = 318 AND Y = 53 else
"000000000000" when X = 319 AND Y = 53 else
"000000000000" when X = 320 AND Y = 53 else
"000000000000" when X = 321 AND Y = 53 else
"000000000000" when X = 322 AND Y = 53 else
"000000000000" when X = 323 AND Y = 53 else
"000000000000" when X = 324 AND Y = 53 else
"100010011101" when X = 0 AND Y = 54 else
"100010011101" when X = 1 AND Y = 54 else
"100010011101" when X = 2 AND Y = 54 else
"100010011101" when X = 3 AND Y = 54 else
"100010011101" when X = 4 AND Y = 54 else
"100010011101" when X = 5 AND Y = 54 else
"100010011101" when X = 6 AND Y = 54 else
"100010011101" when X = 7 AND Y = 54 else
"100010011101" when X = 8 AND Y = 54 else
"100010011101" when X = 9 AND Y = 54 else
"100010011101" when X = 10 AND Y = 54 else
"100010011101" when X = 11 AND Y = 54 else
"100010011101" when X = 12 AND Y = 54 else
"100010011101" when X = 13 AND Y = 54 else
"100010011101" when X = 14 AND Y = 54 else
"100010011101" when X = 15 AND Y = 54 else
"100010011101" when X = 16 AND Y = 54 else
"100010011101" when X = 17 AND Y = 54 else
"100010011101" when X = 18 AND Y = 54 else
"100010011101" when X = 19 AND Y = 54 else
"100010011101" when X = 20 AND Y = 54 else
"100010011101" when X = 21 AND Y = 54 else
"100010011101" when X = 22 AND Y = 54 else
"100010011101" when X = 23 AND Y = 54 else
"100010011101" when X = 24 AND Y = 54 else
"100010011101" when X = 25 AND Y = 54 else
"100010011101" when X = 26 AND Y = 54 else
"100010011101" when X = 27 AND Y = 54 else
"100010011101" when X = 28 AND Y = 54 else
"100010011101" when X = 29 AND Y = 54 else
"100010011101" when X = 30 AND Y = 54 else
"100010011101" when X = 31 AND Y = 54 else
"100010011101" when X = 32 AND Y = 54 else
"100010011101" when X = 33 AND Y = 54 else
"100010011101" when X = 34 AND Y = 54 else
"100010011101" when X = 35 AND Y = 54 else
"100010011101" when X = 36 AND Y = 54 else
"100010011101" when X = 37 AND Y = 54 else
"100010011101" when X = 38 AND Y = 54 else
"100010011101" when X = 39 AND Y = 54 else
"100010011101" when X = 40 AND Y = 54 else
"100010011101" when X = 41 AND Y = 54 else
"100010011101" when X = 42 AND Y = 54 else
"100010011101" when X = 43 AND Y = 54 else
"100010011101" when X = 44 AND Y = 54 else
"110111011111" when X = 45 AND Y = 54 else
"110111011111" when X = 46 AND Y = 54 else
"110111011111" when X = 47 AND Y = 54 else
"110111011111" when X = 48 AND Y = 54 else
"110111011111" when X = 49 AND Y = 54 else
"110111011111" when X = 50 AND Y = 54 else
"110111011111" when X = 51 AND Y = 54 else
"110111011111" when X = 52 AND Y = 54 else
"110111011111" when X = 53 AND Y = 54 else
"110111011111" when X = 54 AND Y = 54 else
"110111011111" when X = 55 AND Y = 54 else
"110111011111" when X = 56 AND Y = 54 else
"110111011111" when X = 57 AND Y = 54 else
"110111011111" when X = 58 AND Y = 54 else
"110111011111" when X = 59 AND Y = 54 else
"110111011111" when X = 60 AND Y = 54 else
"110111011111" when X = 61 AND Y = 54 else
"110111011111" when X = 62 AND Y = 54 else
"110111011111" when X = 63 AND Y = 54 else
"110111011111" when X = 64 AND Y = 54 else
"110111011111" when X = 65 AND Y = 54 else
"110111011111" when X = 66 AND Y = 54 else
"110111011111" when X = 67 AND Y = 54 else
"110111011111" when X = 68 AND Y = 54 else
"110111011111" when X = 69 AND Y = 54 else
"111111111111" when X = 70 AND Y = 54 else
"111111111111" when X = 71 AND Y = 54 else
"111111111111" when X = 72 AND Y = 54 else
"111111111111" when X = 73 AND Y = 54 else
"111111111111" when X = 74 AND Y = 54 else
"111111111111" when X = 75 AND Y = 54 else
"111111111111" when X = 76 AND Y = 54 else
"111111111111" when X = 77 AND Y = 54 else
"111111111111" when X = 78 AND Y = 54 else
"111111111111" when X = 79 AND Y = 54 else
"111111111111" when X = 80 AND Y = 54 else
"111111111111" when X = 81 AND Y = 54 else
"111111111111" when X = 82 AND Y = 54 else
"111111111111" when X = 83 AND Y = 54 else
"111111111111" when X = 84 AND Y = 54 else
"111111111111" when X = 85 AND Y = 54 else
"111111111111" when X = 86 AND Y = 54 else
"111111111111" when X = 87 AND Y = 54 else
"111111111111" when X = 88 AND Y = 54 else
"111111111111" when X = 89 AND Y = 54 else
"111111111111" when X = 90 AND Y = 54 else
"111111111111" when X = 91 AND Y = 54 else
"111111111111" when X = 92 AND Y = 54 else
"111111111111" when X = 93 AND Y = 54 else
"111111111111" when X = 94 AND Y = 54 else
"111111111111" when X = 95 AND Y = 54 else
"111111111111" when X = 96 AND Y = 54 else
"111111111111" when X = 97 AND Y = 54 else
"111111111111" when X = 98 AND Y = 54 else
"111111111111" when X = 99 AND Y = 54 else
"111111111111" when X = 100 AND Y = 54 else
"111111111111" when X = 101 AND Y = 54 else
"111111111111" when X = 102 AND Y = 54 else
"111111111111" when X = 103 AND Y = 54 else
"111111111111" when X = 104 AND Y = 54 else
"111111111111" when X = 105 AND Y = 54 else
"111111111111" when X = 106 AND Y = 54 else
"111111111111" when X = 107 AND Y = 54 else
"111111111111" when X = 108 AND Y = 54 else
"111111111111" when X = 109 AND Y = 54 else
"111111111111" when X = 110 AND Y = 54 else
"111111111111" when X = 111 AND Y = 54 else
"111111111111" when X = 112 AND Y = 54 else
"111111111111" when X = 113 AND Y = 54 else
"111111111111" when X = 114 AND Y = 54 else
"111111111111" when X = 115 AND Y = 54 else
"111111111111" when X = 116 AND Y = 54 else
"111111111111" when X = 117 AND Y = 54 else
"111111111111" when X = 118 AND Y = 54 else
"111111111111" when X = 119 AND Y = 54 else
"111111111111" when X = 120 AND Y = 54 else
"111111111111" when X = 121 AND Y = 54 else
"111111111111" when X = 122 AND Y = 54 else
"111111111111" when X = 123 AND Y = 54 else
"111111111111" when X = 124 AND Y = 54 else
"111111111111" when X = 125 AND Y = 54 else
"111111111111" when X = 126 AND Y = 54 else
"111111111111" when X = 127 AND Y = 54 else
"111111111111" when X = 128 AND Y = 54 else
"111111111111" when X = 129 AND Y = 54 else
"111111111111" when X = 130 AND Y = 54 else
"111111111111" when X = 131 AND Y = 54 else
"111111111111" when X = 132 AND Y = 54 else
"111111111111" when X = 133 AND Y = 54 else
"111111111111" when X = 134 AND Y = 54 else
"111111111111" when X = 135 AND Y = 54 else
"111111111111" when X = 136 AND Y = 54 else
"111111111111" when X = 137 AND Y = 54 else
"111111111111" when X = 138 AND Y = 54 else
"111111111111" when X = 139 AND Y = 54 else
"111111111111" when X = 140 AND Y = 54 else
"111111111111" when X = 141 AND Y = 54 else
"111111111111" when X = 142 AND Y = 54 else
"111111111111" when X = 143 AND Y = 54 else
"111111111111" when X = 144 AND Y = 54 else
"111111111111" when X = 145 AND Y = 54 else
"111111111111" when X = 146 AND Y = 54 else
"111111111111" when X = 147 AND Y = 54 else
"111111111111" when X = 148 AND Y = 54 else
"111111111111" when X = 149 AND Y = 54 else
"111111111111" when X = 150 AND Y = 54 else
"111111111111" when X = 151 AND Y = 54 else
"111111111111" when X = 152 AND Y = 54 else
"111111111111" when X = 153 AND Y = 54 else
"111111111111" when X = 154 AND Y = 54 else
"111111111111" when X = 155 AND Y = 54 else
"111111111111" when X = 156 AND Y = 54 else
"111111111111" when X = 157 AND Y = 54 else
"111111111111" when X = 158 AND Y = 54 else
"111111111111" when X = 159 AND Y = 54 else
"111111111111" when X = 160 AND Y = 54 else
"111111111111" when X = 161 AND Y = 54 else
"111111111111" when X = 162 AND Y = 54 else
"111111111111" when X = 163 AND Y = 54 else
"111111111111" when X = 164 AND Y = 54 else
"111111111111" when X = 165 AND Y = 54 else
"111111111111" when X = 166 AND Y = 54 else
"111111111111" when X = 167 AND Y = 54 else
"111111111111" when X = 168 AND Y = 54 else
"111111111111" when X = 169 AND Y = 54 else
"111111111111" when X = 170 AND Y = 54 else
"111111111111" when X = 171 AND Y = 54 else
"111111111111" when X = 172 AND Y = 54 else
"111111111111" when X = 173 AND Y = 54 else
"111111111111" when X = 174 AND Y = 54 else
"111111111111" when X = 175 AND Y = 54 else
"111111111111" when X = 176 AND Y = 54 else
"111111111111" when X = 177 AND Y = 54 else
"111111111111" when X = 178 AND Y = 54 else
"111111111111" when X = 179 AND Y = 54 else
"111111111111" when X = 180 AND Y = 54 else
"111111111111" when X = 181 AND Y = 54 else
"111111111111" when X = 182 AND Y = 54 else
"111111111111" when X = 183 AND Y = 54 else
"111111111111" when X = 184 AND Y = 54 else
"111111111111" when X = 185 AND Y = 54 else
"111111111111" when X = 186 AND Y = 54 else
"111111111111" when X = 187 AND Y = 54 else
"111111111111" when X = 188 AND Y = 54 else
"111111111111" when X = 189 AND Y = 54 else
"111111111111" when X = 190 AND Y = 54 else
"111111111111" when X = 191 AND Y = 54 else
"111111111111" when X = 192 AND Y = 54 else
"111111111111" when X = 193 AND Y = 54 else
"111111111111" when X = 194 AND Y = 54 else
"111111111111" when X = 195 AND Y = 54 else
"111111111111" when X = 196 AND Y = 54 else
"111111111111" when X = 197 AND Y = 54 else
"111111111111" when X = 198 AND Y = 54 else
"111111111111" when X = 199 AND Y = 54 else
"111111111111" when X = 200 AND Y = 54 else
"111111111111" when X = 201 AND Y = 54 else
"111111111111" when X = 202 AND Y = 54 else
"111111111111" when X = 203 AND Y = 54 else
"111111111111" when X = 204 AND Y = 54 else
"111111111111" when X = 205 AND Y = 54 else
"111111111111" when X = 206 AND Y = 54 else
"111111111111" when X = 207 AND Y = 54 else
"111111111111" when X = 208 AND Y = 54 else
"111111111111" when X = 209 AND Y = 54 else
"111111111111" when X = 210 AND Y = 54 else
"111111111111" when X = 211 AND Y = 54 else
"111111111111" when X = 212 AND Y = 54 else
"111111111111" when X = 213 AND Y = 54 else
"111111111111" when X = 214 AND Y = 54 else
"111111111111" when X = 215 AND Y = 54 else
"111111111111" when X = 216 AND Y = 54 else
"111111111111" when X = 217 AND Y = 54 else
"111111111111" when X = 218 AND Y = 54 else
"111111111111" when X = 219 AND Y = 54 else
"111111111111" when X = 220 AND Y = 54 else
"111111111111" when X = 221 AND Y = 54 else
"111111111111" when X = 222 AND Y = 54 else
"111111111111" when X = 223 AND Y = 54 else
"111111111111" when X = 224 AND Y = 54 else
"111111111111" when X = 225 AND Y = 54 else
"111111111111" when X = 226 AND Y = 54 else
"111111111111" when X = 227 AND Y = 54 else
"111111111111" when X = 228 AND Y = 54 else
"111111111111" when X = 229 AND Y = 54 else
"111111111111" when X = 230 AND Y = 54 else
"111111111111" when X = 231 AND Y = 54 else
"111111111111" when X = 232 AND Y = 54 else
"111111111111" when X = 233 AND Y = 54 else
"111111111111" when X = 234 AND Y = 54 else
"111111111111" when X = 235 AND Y = 54 else
"111111111111" when X = 236 AND Y = 54 else
"111111111111" when X = 237 AND Y = 54 else
"111111111111" when X = 238 AND Y = 54 else
"111111111111" when X = 239 AND Y = 54 else
"111111111111" when X = 240 AND Y = 54 else
"111111111111" when X = 241 AND Y = 54 else
"111111111111" when X = 242 AND Y = 54 else
"111111111111" when X = 243 AND Y = 54 else
"111111111111" when X = 244 AND Y = 54 else
"111111111111" when X = 245 AND Y = 54 else
"111111111111" when X = 246 AND Y = 54 else
"111111111111" when X = 247 AND Y = 54 else
"111111111111" when X = 248 AND Y = 54 else
"111111111111" when X = 249 AND Y = 54 else
"111111111111" when X = 250 AND Y = 54 else
"111111111111" when X = 251 AND Y = 54 else
"111111111111" when X = 252 AND Y = 54 else
"111111111111" when X = 253 AND Y = 54 else
"111111111111" when X = 254 AND Y = 54 else
"111111111111" when X = 255 AND Y = 54 else
"111111111111" when X = 256 AND Y = 54 else
"111111111111" when X = 257 AND Y = 54 else
"111111111111" when X = 258 AND Y = 54 else
"111111111111" when X = 259 AND Y = 54 else
"111111111111" when X = 260 AND Y = 54 else
"111111111111" when X = 261 AND Y = 54 else
"111111111111" when X = 262 AND Y = 54 else
"111111111111" when X = 263 AND Y = 54 else
"111111111111" when X = 264 AND Y = 54 else
"110111011111" when X = 265 AND Y = 54 else
"110111011111" when X = 266 AND Y = 54 else
"110111011111" when X = 267 AND Y = 54 else
"110111011111" when X = 268 AND Y = 54 else
"110111011111" when X = 269 AND Y = 54 else
"110111011111" when X = 270 AND Y = 54 else
"110111011111" when X = 271 AND Y = 54 else
"110111011111" when X = 272 AND Y = 54 else
"110111011111" when X = 273 AND Y = 54 else
"110111011111" when X = 274 AND Y = 54 else
"110111011111" when X = 275 AND Y = 54 else
"110111011111" when X = 276 AND Y = 54 else
"110111011111" when X = 277 AND Y = 54 else
"110111011111" when X = 278 AND Y = 54 else
"110111011111" when X = 279 AND Y = 54 else
"000000000000" when X = 280 AND Y = 54 else
"000000000000" when X = 281 AND Y = 54 else
"000000000000" when X = 282 AND Y = 54 else
"000000000000" when X = 283 AND Y = 54 else
"000000000000" when X = 284 AND Y = 54 else
"000000000000" when X = 285 AND Y = 54 else
"000000000000" when X = 286 AND Y = 54 else
"000000000000" when X = 287 AND Y = 54 else
"000000000000" when X = 288 AND Y = 54 else
"000000000000" when X = 289 AND Y = 54 else
"000000000000" when X = 290 AND Y = 54 else
"000000000000" when X = 291 AND Y = 54 else
"000000000000" when X = 292 AND Y = 54 else
"000000000000" when X = 293 AND Y = 54 else
"000000000000" when X = 294 AND Y = 54 else
"000000000000" when X = 295 AND Y = 54 else
"000000000000" when X = 296 AND Y = 54 else
"000000000000" when X = 297 AND Y = 54 else
"000000000000" when X = 298 AND Y = 54 else
"000000000000" when X = 299 AND Y = 54 else
"000000000000" when X = 300 AND Y = 54 else
"000000000000" when X = 301 AND Y = 54 else
"000000000000" when X = 302 AND Y = 54 else
"000000000000" when X = 303 AND Y = 54 else
"000000000000" when X = 304 AND Y = 54 else
"000000000000" when X = 305 AND Y = 54 else
"000000000000" when X = 306 AND Y = 54 else
"000000000000" when X = 307 AND Y = 54 else
"000000000000" when X = 308 AND Y = 54 else
"000000000000" when X = 309 AND Y = 54 else
"000000000000" when X = 310 AND Y = 54 else
"000000000000" when X = 311 AND Y = 54 else
"000000000000" when X = 312 AND Y = 54 else
"000000000000" when X = 313 AND Y = 54 else
"000000000000" when X = 314 AND Y = 54 else
"000000000000" when X = 315 AND Y = 54 else
"000000000000" when X = 316 AND Y = 54 else
"000000000000" when X = 317 AND Y = 54 else
"000000000000" when X = 318 AND Y = 54 else
"000000000000" when X = 319 AND Y = 54 else
"000000000000" when X = 320 AND Y = 54 else
"000000000000" when X = 321 AND Y = 54 else
"000000000000" when X = 322 AND Y = 54 else
"000000000000" when X = 323 AND Y = 54 else
"000000000000" when X = 324 AND Y = 54 else
"100010011101" when X = 0 AND Y = 55 else
"100010011101" when X = 1 AND Y = 55 else
"100010011101" when X = 2 AND Y = 55 else
"100010011101" when X = 3 AND Y = 55 else
"100010011101" when X = 4 AND Y = 55 else
"100010011101" when X = 5 AND Y = 55 else
"100010011101" when X = 6 AND Y = 55 else
"100010011101" when X = 7 AND Y = 55 else
"100010011101" when X = 8 AND Y = 55 else
"100010011101" when X = 9 AND Y = 55 else
"100010011101" when X = 10 AND Y = 55 else
"100010011101" when X = 11 AND Y = 55 else
"100010011101" when X = 12 AND Y = 55 else
"100010011101" when X = 13 AND Y = 55 else
"100010011101" when X = 14 AND Y = 55 else
"100010011101" when X = 15 AND Y = 55 else
"100010011101" when X = 16 AND Y = 55 else
"100010011101" when X = 17 AND Y = 55 else
"100010011101" when X = 18 AND Y = 55 else
"100010011101" when X = 19 AND Y = 55 else
"100010011101" when X = 20 AND Y = 55 else
"100010011101" when X = 21 AND Y = 55 else
"100010011101" when X = 22 AND Y = 55 else
"100010011101" when X = 23 AND Y = 55 else
"100010011101" when X = 24 AND Y = 55 else
"100010011101" when X = 25 AND Y = 55 else
"100010011101" when X = 26 AND Y = 55 else
"100010011101" when X = 27 AND Y = 55 else
"100010011101" when X = 28 AND Y = 55 else
"100010011101" when X = 29 AND Y = 55 else
"100010011101" when X = 30 AND Y = 55 else
"100010011101" when X = 31 AND Y = 55 else
"100010011101" when X = 32 AND Y = 55 else
"100010011101" when X = 33 AND Y = 55 else
"100010011101" when X = 34 AND Y = 55 else
"100010011101" when X = 35 AND Y = 55 else
"100010011101" when X = 36 AND Y = 55 else
"100010011101" when X = 37 AND Y = 55 else
"100010011101" when X = 38 AND Y = 55 else
"100010011101" when X = 39 AND Y = 55 else
"110111011111" when X = 40 AND Y = 55 else
"110111011111" when X = 41 AND Y = 55 else
"110111011111" when X = 42 AND Y = 55 else
"110111011111" when X = 43 AND Y = 55 else
"110111011111" when X = 44 AND Y = 55 else
"110111011111" when X = 45 AND Y = 55 else
"110111011111" when X = 46 AND Y = 55 else
"110111011111" when X = 47 AND Y = 55 else
"110111011111" when X = 48 AND Y = 55 else
"110111011111" when X = 49 AND Y = 55 else
"110111011111" when X = 50 AND Y = 55 else
"110111011111" when X = 51 AND Y = 55 else
"110111011111" when X = 52 AND Y = 55 else
"110111011111" when X = 53 AND Y = 55 else
"110111011111" when X = 54 AND Y = 55 else
"110111011111" when X = 55 AND Y = 55 else
"110111011111" when X = 56 AND Y = 55 else
"110111011111" when X = 57 AND Y = 55 else
"110111011111" when X = 58 AND Y = 55 else
"110111011111" when X = 59 AND Y = 55 else
"110111011111" when X = 60 AND Y = 55 else
"110111011111" when X = 61 AND Y = 55 else
"110111011111" when X = 62 AND Y = 55 else
"110111011111" when X = 63 AND Y = 55 else
"110111011111" when X = 64 AND Y = 55 else
"110111011111" when X = 65 AND Y = 55 else
"110111011111" when X = 66 AND Y = 55 else
"110111011111" when X = 67 AND Y = 55 else
"110111011111" when X = 68 AND Y = 55 else
"110111011111" when X = 69 AND Y = 55 else
"110111011111" when X = 70 AND Y = 55 else
"110111011111" when X = 71 AND Y = 55 else
"110111011111" when X = 72 AND Y = 55 else
"110111011111" when X = 73 AND Y = 55 else
"110111011111" when X = 74 AND Y = 55 else
"110111011111" when X = 75 AND Y = 55 else
"110111011111" when X = 76 AND Y = 55 else
"110111011111" when X = 77 AND Y = 55 else
"110111011111" when X = 78 AND Y = 55 else
"110111011111" when X = 79 AND Y = 55 else
"110111011111" when X = 80 AND Y = 55 else
"110111011111" when X = 81 AND Y = 55 else
"110111011111" when X = 82 AND Y = 55 else
"110111011111" when X = 83 AND Y = 55 else
"110111011111" when X = 84 AND Y = 55 else
"110111011111" when X = 85 AND Y = 55 else
"110111011111" when X = 86 AND Y = 55 else
"110111011111" when X = 87 AND Y = 55 else
"110111011111" when X = 88 AND Y = 55 else
"110111011111" when X = 89 AND Y = 55 else
"110111011111" when X = 90 AND Y = 55 else
"110111011111" when X = 91 AND Y = 55 else
"110111011111" when X = 92 AND Y = 55 else
"110111011111" when X = 93 AND Y = 55 else
"110111011111" when X = 94 AND Y = 55 else
"111111111111" when X = 95 AND Y = 55 else
"111111111111" when X = 96 AND Y = 55 else
"111111111111" when X = 97 AND Y = 55 else
"111111111111" when X = 98 AND Y = 55 else
"111111111111" when X = 99 AND Y = 55 else
"111111111111" when X = 100 AND Y = 55 else
"111111111111" when X = 101 AND Y = 55 else
"111111111111" when X = 102 AND Y = 55 else
"111111111111" when X = 103 AND Y = 55 else
"111111111111" when X = 104 AND Y = 55 else
"111111111111" when X = 105 AND Y = 55 else
"111111111111" when X = 106 AND Y = 55 else
"111111111111" when X = 107 AND Y = 55 else
"111111111111" when X = 108 AND Y = 55 else
"111111111111" when X = 109 AND Y = 55 else
"111111111111" when X = 110 AND Y = 55 else
"111111111111" when X = 111 AND Y = 55 else
"111111111111" when X = 112 AND Y = 55 else
"111111111111" when X = 113 AND Y = 55 else
"111111111111" when X = 114 AND Y = 55 else
"111111111111" when X = 115 AND Y = 55 else
"111111111111" when X = 116 AND Y = 55 else
"111111111111" when X = 117 AND Y = 55 else
"111111111111" when X = 118 AND Y = 55 else
"111111111111" when X = 119 AND Y = 55 else
"111111111111" when X = 120 AND Y = 55 else
"111111111111" when X = 121 AND Y = 55 else
"111111111111" when X = 122 AND Y = 55 else
"111111111111" when X = 123 AND Y = 55 else
"111111111111" when X = 124 AND Y = 55 else
"111111111111" when X = 125 AND Y = 55 else
"111111111111" when X = 126 AND Y = 55 else
"111111111111" when X = 127 AND Y = 55 else
"111111111111" when X = 128 AND Y = 55 else
"111111111111" when X = 129 AND Y = 55 else
"111111111111" when X = 130 AND Y = 55 else
"111111111111" when X = 131 AND Y = 55 else
"111111111111" when X = 132 AND Y = 55 else
"111111111111" when X = 133 AND Y = 55 else
"111111111111" when X = 134 AND Y = 55 else
"111111111111" when X = 135 AND Y = 55 else
"111111111111" when X = 136 AND Y = 55 else
"111111111111" when X = 137 AND Y = 55 else
"111111111111" when X = 138 AND Y = 55 else
"111111111111" when X = 139 AND Y = 55 else
"111111111111" when X = 140 AND Y = 55 else
"111111111111" when X = 141 AND Y = 55 else
"111111111111" when X = 142 AND Y = 55 else
"111111111111" when X = 143 AND Y = 55 else
"111111111111" when X = 144 AND Y = 55 else
"111111111111" when X = 145 AND Y = 55 else
"111111111111" when X = 146 AND Y = 55 else
"111111111111" when X = 147 AND Y = 55 else
"111111111111" when X = 148 AND Y = 55 else
"111111111111" when X = 149 AND Y = 55 else
"111111111111" when X = 150 AND Y = 55 else
"111111111111" when X = 151 AND Y = 55 else
"111111111111" when X = 152 AND Y = 55 else
"111111111111" when X = 153 AND Y = 55 else
"111111111111" when X = 154 AND Y = 55 else
"111111111111" when X = 155 AND Y = 55 else
"111111111111" when X = 156 AND Y = 55 else
"111111111111" when X = 157 AND Y = 55 else
"111111111111" when X = 158 AND Y = 55 else
"111111111111" when X = 159 AND Y = 55 else
"111111111111" when X = 160 AND Y = 55 else
"111111111111" when X = 161 AND Y = 55 else
"111111111111" when X = 162 AND Y = 55 else
"111111111111" when X = 163 AND Y = 55 else
"111111111111" when X = 164 AND Y = 55 else
"111111111111" when X = 165 AND Y = 55 else
"111111111111" when X = 166 AND Y = 55 else
"111111111111" when X = 167 AND Y = 55 else
"111111111111" when X = 168 AND Y = 55 else
"111111111111" when X = 169 AND Y = 55 else
"111111111111" when X = 170 AND Y = 55 else
"111111111111" when X = 171 AND Y = 55 else
"111111111111" when X = 172 AND Y = 55 else
"111111111111" when X = 173 AND Y = 55 else
"111111111111" when X = 174 AND Y = 55 else
"111111111111" when X = 175 AND Y = 55 else
"111111111111" when X = 176 AND Y = 55 else
"111111111111" when X = 177 AND Y = 55 else
"111111111111" when X = 178 AND Y = 55 else
"111111111111" when X = 179 AND Y = 55 else
"111111111111" when X = 180 AND Y = 55 else
"111111111111" when X = 181 AND Y = 55 else
"111111111111" when X = 182 AND Y = 55 else
"111111111111" when X = 183 AND Y = 55 else
"111111111111" when X = 184 AND Y = 55 else
"111111111111" when X = 185 AND Y = 55 else
"111111111111" when X = 186 AND Y = 55 else
"111111111111" when X = 187 AND Y = 55 else
"111111111111" when X = 188 AND Y = 55 else
"111111111111" when X = 189 AND Y = 55 else
"111111111111" when X = 190 AND Y = 55 else
"111111111111" when X = 191 AND Y = 55 else
"111111111111" when X = 192 AND Y = 55 else
"111111111111" when X = 193 AND Y = 55 else
"111111111111" when X = 194 AND Y = 55 else
"111111111111" when X = 195 AND Y = 55 else
"111111111111" when X = 196 AND Y = 55 else
"111111111111" when X = 197 AND Y = 55 else
"111111111111" when X = 198 AND Y = 55 else
"111111111111" when X = 199 AND Y = 55 else
"111111111111" when X = 200 AND Y = 55 else
"111111111111" when X = 201 AND Y = 55 else
"111111111111" when X = 202 AND Y = 55 else
"111111111111" when X = 203 AND Y = 55 else
"111111111111" when X = 204 AND Y = 55 else
"111111111111" when X = 205 AND Y = 55 else
"111111111111" when X = 206 AND Y = 55 else
"111111111111" when X = 207 AND Y = 55 else
"111111111111" when X = 208 AND Y = 55 else
"111111111111" when X = 209 AND Y = 55 else
"111111111111" when X = 210 AND Y = 55 else
"111111111111" when X = 211 AND Y = 55 else
"111111111111" when X = 212 AND Y = 55 else
"111111111111" when X = 213 AND Y = 55 else
"111111111111" when X = 214 AND Y = 55 else
"111111111111" when X = 215 AND Y = 55 else
"111111111111" when X = 216 AND Y = 55 else
"111111111111" when X = 217 AND Y = 55 else
"111111111111" when X = 218 AND Y = 55 else
"111111111111" when X = 219 AND Y = 55 else
"111111111111" when X = 220 AND Y = 55 else
"111111111111" when X = 221 AND Y = 55 else
"111111111111" when X = 222 AND Y = 55 else
"111111111111" when X = 223 AND Y = 55 else
"111111111111" when X = 224 AND Y = 55 else
"111111111111" when X = 225 AND Y = 55 else
"111111111111" when X = 226 AND Y = 55 else
"111111111111" when X = 227 AND Y = 55 else
"111111111111" when X = 228 AND Y = 55 else
"111111111111" when X = 229 AND Y = 55 else
"111111111111" when X = 230 AND Y = 55 else
"111111111111" when X = 231 AND Y = 55 else
"111111111111" when X = 232 AND Y = 55 else
"111111111111" when X = 233 AND Y = 55 else
"111111111111" when X = 234 AND Y = 55 else
"111111111111" when X = 235 AND Y = 55 else
"111111111111" when X = 236 AND Y = 55 else
"111111111111" when X = 237 AND Y = 55 else
"111111111111" when X = 238 AND Y = 55 else
"111111111111" when X = 239 AND Y = 55 else
"111111111111" when X = 240 AND Y = 55 else
"111111111111" when X = 241 AND Y = 55 else
"111111111111" when X = 242 AND Y = 55 else
"111111111111" when X = 243 AND Y = 55 else
"111111111111" when X = 244 AND Y = 55 else
"111111111111" when X = 245 AND Y = 55 else
"111111111111" when X = 246 AND Y = 55 else
"111111111111" when X = 247 AND Y = 55 else
"111111111111" when X = 248 AND Y = 55 else
"111111111111" when X = 249 AND Y = 55 else
"111111111111" when X = 250 AND Y = 55 else
"111111111111" when X = 251 AND Y = 55 else
"111111111111" when X = 252 AND Y = 55 else
"111111111111" when X = 253 AND Y = 55 else
"111111111111" when X = 254 AND Y = 55 else
"111111111111" when X = 255 AND Y = 55 else
"111111111111" when X = 256 AND Y = 55 else
"111111111111" when X = 257 AND Y = 55 else
"111111111111" when X = 258 AND Y = 55 else
"111111111111" when X = 259 AND Y = 55 else
"111111111111" when X = 260 AND Y = 55 else
"111111111111" when X = 261 AND Y = 55 else
"111111111111" when X = 262 AND Y = 55 else
"111111111111" when X = 263 AND Y = 55 else
"111111111111" when X = 264 AND Y = 55 else
"110111011111" when X = 265 AND Y = 55 else
"110111011111" when X = 266 AND Y = 55 else
"110111011111" when X = 267 AND Y = 55 else
"110111011111" when X = 268 AND Y = 55 else
"110111011111" when X = 269 AND Y = 55 else
"110111011111" when X = 270 AND Y = 55 else
"110111011111" when X = 271 AND Y = 55 else
"110111011111" when X = 272 AND Y = 55 else
"110111011111" when X = 273 AND Y = 55 else
"110111011111" when X = 274 AND Y = 55 else
"110111011111" when X = 275 AND Y = 55 else
"110111011111" when X = 276 AND Y = 55 else
"110111011111" when X = 277 AND Y = 55 else
"110111011111" when X = 278 AND Y = 55 else
"110111011111" when X = 279 AND Y = 55 else
"000000000000" when X = 280 AND Y = 55 else
"000000000000" when X = 281 AND Y = 55 else
"000000000000" when X = 282 AND Y = 55 else
"000000000000" when X = 283 AND Y = 55 else
"000000000000" when X = 284 AND Y = 55 else
"000000000000" when X = 285 AND Y = 55 else
"000000000000" when X = 286 AND Y = 55 else
"000000000000" when X = 287 AND Y = 55 else
"000000000000" when X = 288 AND Y = 55 else
"000000000000" when X = 289 AND Y = 55 else
"000000000000" when X = 290 AND Y = 55 else
"000000000000" when X = 291 AND Y = 55 else
"000000000000" when X = 292 AND Y = 55 else
"000000000000" when X = 293 AND Y = 55 else
"000000000000" when X = 294 AND Y = 55 else
"000000000000" when X = 295 AND Y = 55 else
"000000000000" when X = 296 AND Y = 55 else
"000000000000" when X = 297 AND Y = 55 else
"000000000000" when X = 298 AND Y = 55 else
"000000000000" when X = 299 AND Y = 55 else
"000000000000" when X = 300 AND Y = 55 else
"000000000000" when X = 301 AND Y = 55 else
"000000000000" when X = 302 AND Y = 55 else
"000000000000" when X = 303 AND Y = 55 else
"000000000000" when X = 304 AND Y = 55 else
"000000000000" when X = 305 AND Y = 55 else
"000000000000" when X = 306 AND Y = 55 else
"000000000000" when X = 307 AND Y = 55 else
"000000000000" when X = 308 AND Y = 55 else
"000000000000" when X = 309 AND Y = 55 else
"000000000000" when X = 310 AND Y = 55 else
"000000000000" when X = 311 AND Y = 55 else
"000000000000" when X = 312 AND Y = 55 else
"000000000000" when X = 313 AND Y = 55 else
"000000000000" when X = 314 AND Y = 55 else
"000000000000" when X = 315 AND Y = 55 else
"000000000000" when X = 316 AND Y = 55 else
"000000000000" when X = 317 AND Y = 55 else
"000000000000" when X = 318 AND Y = 55 else
"000000000000" when X = 319 AND Y = 55 else
"000000000000" when X = 320 AND Y = 55 else
"000000000000" when X = 321 AND Y = 55 else
"000000000000" when X = 322 AND Y = 55 else
"000000000000" when X = 323 AND Y = 55 else
"000000000000" when X = 324 AND Y = 55 else
"100010011101" when X = 0 AND Y = 56 else
"100010011101" when X = 1 AND Y = 56 else
"100010011101" when X = 2 AND Y = 56 else
"100010011101" when X = 3 AND Y = 56 else
"100010011101" when X = 4 AND Y = 56 else
"100010011101" when X = 5 AND Y = 56 else
"100010011101" when X = 6 AND Y = 56 else
"100010011101" when X = 7 AND Y = 56 else
"100010011101" when X = 8 AND Y = 56 else
"100010011101" when X = 9 AND Y = 56 else
"100010011101" when X = 10 AND Y = 56 else
"100010011101" when X = 11 AND Y = 56 else
"100010011101" when X = 12 AND Y = 56 else
"100010011101" when X = 13 AND Y = 56 else
"100010011101" when X = 14 AND Y = 56 else
"100010011101" when X = 15 AND Y = 56 else
"100010011101" when X = 16 AND Y = 56 else
"100010011101" when X = 17 AND Y = 56 else
"100010011101" when X = 18 AND Y = 56 else
"100010011101" when X = 19 AND Y = 56 else
"100010011101" when X = 20 AND Y = 56 else
"100010011101" when X = 21 AND Y = 56 else
"100010011101" when X = 22 AND Y = 56 else
"100010011101" when X = 23 AND Y = 56 else
"100010011101" when X = 24 AND Y = 56 else
"100010011101" when X = 25 AND Y = 56 else
"100010011101" when X = 26 AND Y = 56 else
"100010011101" when X = 27 AND Y = 56 else
"100010011101" when X = 28 AND Y = 56 else
"100010011101" when X = 29 AND Y = 56 else
"100010011101" when X = 30 AND Y = 56 else
"100010011101" when X = 31 AND Y = 56 else
"100010011101" when X = 32 AND Y = 56 else
"100010011101" when X = 33 AND Y = 56 else
"100010011101" when X = 34 AND Y = 56 else
"100010011101" when X = 35 AND Y = 56 else
"100010011101" when X = 36 AND Y = 56 else
"100010011101" when X = 37 AND Y = 56 else
"100010011101" when X = 38 AND Y = 56 else
"100010011101" when X = 39 AND Y = 56 else
"110111011111" when X = 40 AND Y = 56 else
"110111011111" when X = 41 AND Y = 56 else
"110111011111" when X = 42 AND Y = 56 else
"110111011111" when X = 43 AND Y = 56 else
"110111011111" when X = 44 AND Y = 56 else
"110111011111" when X = 45 AND Y = 56 else
"110111011111" when X = 46 AND Y = 56 else
"110111011111" when X = 47 AND Y = 56 else
"110111011111" when X = 48 AND Y = 56 else
"110111011111" when X = 49 AND Y = 56 else
"110111011111" when X = 50 AND Y = 56 else
"110111011111" when X = 51 AND Y = 56 else
"110111011111" when X = 52 AND Y = 56 else
"110111011111" when X = 53 AND Y = 56 else
"110111011111" when X = 54 AND Y = 56 else
"110111011111" when X = 55 AND Y = 56 else
"110111011111" when X = 56 AND Y = 56 else
"110111011111" when X = 57 AND Y = 56 else
"110111011111" when X = 58 AND Y = 56 else
"110111011111" when X = 59 AND Y = 56 else
"110111011111" when X = 60 AND Y = 56 else
"110111011111" when X = 61 AND Y = 56 else
"110111011111" when X = 62 AND Y = 56 else
"110111011111" when X = 63 AND Y = 56 else
"110111011111" when X = 64 AND Y = 56 else
"110111011111" when X = 65 AND Y = 56 else
"110111011111" when X = 66 AND Y = 56 else
"110111011111" when X = 67 AND Y = 56 else
"110111011111" when X = 68 AND Y = 56 else
"110111011111" when X = 69 AND Y = 56 else
"110111011111" when X = 70 AND Y = 56 else
"110111011111" when X = 71 AND Y = 56 else
"110111011111" when X = 72 AND Y = 56 else
"110111011111" when X = 73 AND Y = 56 else
"110111011111" when X = 74 AND Y = 56 else
"110111011111" when X = 75 AND Y = 56 else
"110111011111" when X = 76 AND Y = 56 else
"110111011111" when X = 77 AND Y = 56 else
"110111011111" when X = 78 AND Y = 56 else
"110111011111" when X = 79 AND Y = 56 else
"110111011111" when X = 80 AND Y = 56 else
"110111011111" when X = 81 AND Y = 56 else
"110111011111" when X = 82 AND Y = 56 else
"110111011111" when X = 83 AND Y = 56 else
"110111011111" when X = 84 AND Y = 56 else
"110111011111" when X = 85 AND Y = 56 else
"110111011111" when X = 86 AND Y = 56 else
"110111011111" when X = 87 AND Y = 56 else
"110111011111" when X = 88 AND Y = 56 else
"110111011111" when X = 89 AND Y = 56 else
"110111011111" when X = 90 AND Y = 56 else
"110111011111" when X = 91 AND Y = 56 else
"110111011111" when X = 92 AND Y = 56 else
"110111011111" when X = 93 AND Y = 56 else
"110111011111" when X = 94 AND Y = 56 else
"111111111111" when X = 95 AND Y = 56 else
"111111111111" when X = 96 AND Y = 56 else
"111111111111" when X = 97 AND Y = 56 else
"111111111111" when X = 98 AND Y = 56 else
"111111111111" when X = 99 AND Y = 56 else
"111111111111" when X = 100 AND Y = 56 else
"111111111111" when X = 101 AND Y = 56 else
"111111111111" when X = 102 AND Y = 56 else
"111111111111" when X = 103 AND Y = 56 else
"111111111111" when X = 104 AND Y = 56 else
"111111111111" when X = 105 AND Y = 56 else
"111111111111" when X = 106 AND Y = 56 else
"111111111111" when X = 107 AND Y = 56 else
"111111111111" when X = 108 AND Y = 56 else
"111111111111" when X = 109 AND Y = 56 else
"111111111111" when X = 110 AND Y = 56 else
"111111111111" when X = 111 AND Y = 56 else
"111111111111" when X = 112 AND Y = 56 else
"111111111111" when X = 113 AND Y = 56 else
"111111111111" when X = 114 AND Y = 56 else
"111111111111" when X = 115 AND Y = 56 else
"111111111111" when X = 116 AND Y = 56 else
"111111111111" when X = 117 AND Y = 56 else
"111111111111" when X = 118 AND Y = 56 else
"111111111111" when X = 119 AND Y = 56 else
"111111111111" when X = 120 AND Y = 56 else
"111111111111" when X = 121 AND Y = 56 else
"111111111111" when X = 122 AND Y = 56 else
"111111111111" when X = 123 AND Y = 56 else
"111111111111" when X = 124 AND Y = 56 else
"111111111111" when X = 125 AND Y = 56 else
"111111111111" when X = 126 AND Y = 56 else
"111111111111" when X = 127 AND Y = 56 else
"111111111111" when X = 128 AND Y = 56 else
"111111111111" when X = 129 AND Y = 56 else
"111111111111" when X = 130 AND Y = 56 else
"111111111111" when X = 131 AND Y = 56 else
"111111111111" when X = 132 AND Y = 56 else
"111111111111" when X = 133 AND Y = 56 else
"111111111111" when X = 134 AND Y = 56 else
"111111111111" when X = 135 AND Y = 56 else
"111111111111" when X = 136 AND Y = 56 else
"111111111111" when X = 137 AND Y = 56 else
"111111111111" when X = 138 AND Y = 56 else
"111111111111" when X = 139 AND Y = 56 else
"111111111111" when X = 140 AND Y = 56 else
"111111111111" when X = 141 AND Y = 56 else
"111111111111" when X = 142 AND Y = 56 else
"111111111111" when X = 143 AND Y = 56 else
"111111111111" when X = 144 AND Y = 56 else
"111111111111" when X = 145 AND Y = 56 else
"111111111111" when X = 146 AND Y = 56 else
"111111111111" when X = 147 AND Y = 56 else
"111111111111" when X = 148 AND Y = 56 else
"111111111111" when X = 149 AND Y = 56 else
"111111111111" when X = 150 AND Y = 56 else
"111111111111" when X = 151 AND Y = 56 else
"111111111111" when X = 152 AND Y = 56 else
"111111111111" when X = 153 AND Y = 56 else
"111111111111" when X = 154 AND Y = 56 else
"111111111111" when X = 155 AND Y = 56 else
"111111111111" when X = 156 AND Y = 56 else
"111111111111" when X = 157 AND Y = 56 else
"111111111111" when X = 158 AND Y = 56 else
"111111111111" when X = 159 AND Y = 56 else
"111111111111" when X = 160 AND Y = 56 else
"111111111111" when X = 161 AND Y = 56 else
"111111111111" when X = 162 AND Y = 56 else
"111111111111" when X = 163 AND Y = 56 else
"111111111111" when X = 164 AND Y = 56 else
"111111111111" when X = 165 AND Y = 56 else
"111111111111" when X = 166 AND Y = 56 else
"111111111111" when X = 167 AND Y = 56 else
"111111111111" when X = 168 AND Y = 56 else
"111111111111" when X = 169 AND Y = 56 else
"111111111111" when X = 170 AND Y = 56 else
"111111111111" when X = 171 AND Y = 56 else
"111111111111" when X = 172 AND Y = 56 else
"111111111111" when X = 173 AND Y = 56 else
"111111111111" when X = 174 AND Y = 56 else
"111111111111" when X = 175 AND Y = 56 else
"111111111111" when X = 176 AND Y = 56 else
"111111111111" when X = 177 AND Y = 56 else
"111111111111" when X = 178 AND Y = 56 else
"111111111111" when X = 179 AND Y = 56 else
"111111111111" when X = 180 AND Y = 56 else
"111111111111" when X = 181 AND Y = 56 else
"111111111111" when X = 182 AND Y = 56 else
"111111111111" when X = 183 AND Y = 56 else
"111111111111" when X = 184 AND Y = 56 else
"111111111111" when X = 185 AND Y = 56 else
"111111111111" when X = 186 AND Y = 56 else
"111111111111" when X = 187 AND Y = 56 else
"111111111111" when X = 188 AND Y = 56 else
"111111111111" when X = 189 AND Y = 56 else
"111111111111" when X = 190 AND Y = 56 else
"111111111111" when X = 191 AND Y = 56 else
"111111111111" when X = 192 AND Y = 56 else
"111111111111" when X = 193 AND Y = 56 else
"111111111111" when X = 194 AND Y = 56 else
"111111111111" when X = 195 AND Y = 56 else
"111111111111" when X = 196 AND Y = 56 else
"111111111111" when X = 197 AND Y = 56 else
"111111111111" when X = 198 AND Y = 56 else
"111111111111" when X = 199 AND Y = 56 else
"111111111111" when X = 200 AND Y = 56 else
"111111111111" when X = 201 AND Y = 56 else
"111111111111" when X = 202 AND Y = 56 else
"111111111111" when X = 203 AND Y = 56 else
"111111111111" when X = 204 AND Y = 56 else
"111111111111" when X = 205 AND Y = 56 else
"111111111111" when X = 206 AND Y = 56 else
"111111111111" when X = 207 AND Y = 56 else
"111111111111" when X = 208 AND Y = 56 else
"111111111111" when X = 209 AND Y = 56 else
"111111111111" when X = 210 AND Y = 56 else
"111111111111" when X = 211 AND Y = 56 else
"111111111111" when X = 212 AND Y = 56 else
"111111111111" when X = 213 AND Y = 56 else
"111111111111" when X = 214 AND Y = 56 else
"111111111111" when X = 215 AND Y = 56 else
"111111111111" when X = 216 AND Y = 56 else
"111111111111" when X = 217 AND Y = 56 else
"111111111111" when X = 218 AND Y = 56 else
"111111111111" when X = 219 AND Y = 56 else
"111111111111" when X = 220 AND Y = 56 else
"111111111111" when X = 221 AND Y = 56 else
"111111111111" when X = 222 AND Y = 56 else
"111111111111" when X = 223 AND Y = 56 else
"111111111111" when X = 224 AND Y = 56 else
"111111111111" when X = 225 AND Y = 56 else
"111111111111" when X = 226 AND Y = 56 else
"111111111111" when X = 227 AND Y = 56 else
"111111111111" when X = 228 AND Y = 56 else
"111111111111" when X = 229 AND Y = 56 else
"111111111111" when X = 230 AND Y = 56 else
"111111111111" when X = 231 AND Y = 56 else
"111111111111" when X = 232 AND Y = 56 else
"111111111111" when X = 233 AND Y = 56 else
"111111111111" when X = 234 AND Y = 56 else
"111111111111" when X = 235 AND Y = 56 else
"111111111111" when X = 236 AND Y = 56 else
"111111111111" when X = 237 AND Y = 56 else
"111111111111" when X = 238 AND Y = 56 else
"111111111111" when X = 239 AND Y = 56 else
"111111111111" when X = 240 AND Y = 56 else
"111111111111" when X = 241 AND Y = 56 else
"111111111111" when X = 242 AND Y = 56 else
"111111111111" when X = 243 AND Y = 56 else
"111111111111" when X = 244 AND Y = 56 else
"111111111111" when X = 245 AND Y = 56 else
"111111111111" when X = 246 AND Y = 56 else
"111111111111" when X = 247 AND Y = 56 else
"111111111111" when X = 248 AND Y = 56 else
"111111111111" when X = 249 AND Y = 56 else
"111111111111" when X = 250 AND Y = 56 else
"111111111111" when X = 251 AND Y = 56 else
"111111111111" when X = 252 AND Y = 56 else
"111111111111" when X = 253 AND Y = 56 else
"111111111111" when X = 254 AND Y = 56 else
"111111111111" when X = 255 AND Y = 56 else
"111111111111" when X = 256 AND Y = 56 else
"111111111111" when X = 257 AND Y = 56 else
"111111111111" when X = 258 AND Y = 56 else
"111111111111" when X = 259 AND Y = 56 else
"111111111111" when X = 260 AND Y = 56 else
"111111111111" when X = 261 AND Y = 56 else
"111111111111" when X = 262 AND Y = 56 else
"111111111111" when X = 263 AND Y = 56 else
"111111111111" when X = 264 AND Y = 56 else
"110111011111" when X = 265 AND Y = 56 else
"110111011111" when X = 266 AND Y = 56 else
"110111011111" when X = 267 AND Y = 56 else
"110111011111" when X = 268 AND Y = 56 else
"110111011111" when X = 269 AND Y = 56 else
"110111011111" when X = 270 AND Y = 56 else
"110111011111" when X = 271 AND Y = 56 else
"110111011111" when X = 272 AND Y = 56 else
"110111011111" when X = 273 AND Y = 56 else
"110111011111" when X = 274 AND Y = 56 else
"110111011111" when X = 275 AND Y = 56 else
"110111011111" when X = 276 AND Y = 56 else
"110111011111" when X = 277 AND Y = 56 else
"110111011111" when X = 278 AND Y = 56 else
"110111011111" when X = 279 AND Y = 56 else
"000000000000" when X = 280 AND Y = 56 else
"000000000000" when X = 281 AND Y = 56 else
"000000000000" when X = 282 AND Y = 56 else
"000000000000" when X = 283 AND Y = 56 else
"000000000000" when X = 284 AND Y = 56 else
"000000000000" when X = 285 AND Y = 56 else
"000000000000" when X = 286 AND Y = 56 else
"000000000000" when X = 287 AND Y = 56 else
"000000000000" when X = 288 AND Y = 56 else
"000000000000" when X = 289 AND Y = 56 else
"000000000000" when X = 290 AND Y = 56 else
"000000000000" when X = 291 AND Y = 56 else
"000000000000" when X = 292 AND Y = 56 else
"000000000000" when X = 293 AND Y = 56 else
"000000000000" when X = 294 AND Y = 56 else
"000000000000" when X = 295 AND Y = 56 else
"000000000000" when X = 296 AND Y = 56 else
"000000000000" when X = 297 AND Y = 56 else
"000000000000" when X = 298 AND Y = 56 else
"000000000000" when X = 299 AND Y = 56 else
"000000000000" when X = 300 AND Y = 56 else
"000000000000" when X = 301 AND Y = 56 else
"000000000000" when X = 302 AND Y = 56 else
"000000000000" when X = 303 AND Y = 56 else
"000000000000" when X = 304 AND Y = 56 else
"000000000000" when X = 305 AND Y = 56 else
"000000000000" when X = 306 AND Y = 56 else
"000000000000" when X = 307 AND Y = 56 else
"000000000000" when X = 308 AND Y = 56 else
"000000000000" when X = 309 AND Y = 56 else
"000000000000" when X = 310 AND Y = 56 else
"000000000000" when X = 311 AND Y = 56 else
"000000000000" when X = 312 AND Y = 56 else
"000000000000" when X = 313 AND Y = 56 else
"000000000000" when X = 314 AND Y = 56 else
"000000000000" when X = 315 AND Y = 56 else
"000000000000" when X = 316 AND Y = 56 else
"000000000000" when X = 317 AND Y = 56 else
"000000000000" when X = 318 AND Y = 56 else
"000000000000" when X = 319 AND Y = 56 else
"000000000000" when X = 320 AND Y = 56 else
"000000000000" when X = 321 AND Y = 56 else
"000000000000" when X = 322 AND Y = 56 else
"000000000000" when X = 323 AND Y = 56 else
"000000000000" when X = 324 AND Y = 56 else
"100010011101" when X = 0 AND Y = 57 else
"100010011101" when X = 1 AND Y = 57 else
"100010011101" when X = 2 AND Y = 57 else
"100010011101" when X = 3 AND Y = 57 else
"100010011101" when X = 4 AND Y = 57 else
"100010011101" when X = 5 AND Y = 57 else
"100010011101" when X = 6 AND Y = 57 else
"100010011101" when X = 7 AND Y = 57 else
"100010011101" when X = 8 AND Y = 57 else
"100010011101" when X = 9 AND Y = 57 else
"100010011101" when X = 10 AND Y = 57 else
"100010011101" when X = 11 AND Y = 57 else
"100010011101" when X = 12 AND Y = 57 else
"100010011101" when X = 13 AND Y = 57 else
"100010011101" when X = 14 AND Y = 57 else
"100010011101" when X = 15 AND Y = 57 else
"100010011101" when X = 16 AND Y = 57 else
"100010011101" when X = 17 AND Y = 57 else
"100010011101" when X = 18 AND Y = 57 else
"100010011101" when X = 19 AND Y = 57 else
"100010011101" when X = 20 AND Y = 57 else
"100010011101" when X = 21 AND Y = 57 else
"100010011101" when X = 22 AND Y = 57 else
"100010011101" when X = 23 AND Y = 57 else
"100010011101" when X = 24 AND Y = 57 else
"100010011101" when X = 25 AND Y = 57 else
"100010011101" when X = 26 AND Y = 57 else
"100010011101" when X = 27 AND Y = 57 else
"100010011101" when X = 28 AND Y = 57 else
"100010011101" when X = 29 AND Y = 57 else
"100010011101" when X = 30 AND Y = 57 else
"100010011101" when X = 31 AND Y = 57 else
"100010011101" when X = 32 AND Y = 57 else
"100010011101" when X = 33 AND Y = 57 else
"100010011101" when X = 34 AND Y = 57 else
"100010011101" when X = 35 AND Y = 57 else
"100010011101" when X = 36 AND Y = 57 else
"100010011101" when X = 37 AND Y = 57 else
"100010011101" when X = 38 AND Y = 57 else
"100010011101" when X = 39 AND Y = 57 else
"110111011111" when X = 40 AND Y = 57 else
"110111011111" when X = 41 AND Y = 57 else
"110111011111" when X = 42 AND Y = 57 else
"110111011111" when X = 43 AND Y = 57 else
"110111011111" when X = 44 AND Y = 57 else
"110111011111" when X = 45 AND Y = 57 else
"110111011111" when X = 46 AND Y = 57 else
"110111011111" when X = 47 AND Y = 57 else
"110111011111" when X = 48 AND Y = 57 else
"110111011111" when X = 49 AND Y = 57 else
"110111011111" when X = 50 AND Y = 57 else
"110111011111" when X = 51 AND Y = 57 else
"110111011111" when X = 52 AND Y = 57 else
"110111011111" when X = 53 AND Y = 57 else
"110111011111" when X = 54 AND Y = 57 else
"110111011111" when X = 55 AND Y = 57 else
"110111011111" when X = 56 AND Y = 57 else
"110111011111" when X = 57 AND Y = 57 else
"110111011111" when X = 58 AND Y = 57 else
"110111011111" when X = 59 AND Y = 57 else
"110111011111" when X = 60 AND Y = 57 else
"110111011111" when X = 61 AND Y = 57 else
"110111011111" when X = 62 AND Y = 57 else
"110111011111" when X = 63 AND Y = 57 else
"110111011111" when X = 64 AND Y = 57 else
"110111011111" when X = 65 AND Y = 57 else
"110111011111" when X = 66 AND Y = 57 else
"110111011111" when X = 67 AND Y = 57 else
"110111011111" when X = 68 AND Y = 57 else
"110111011111" when X = 69 AND Y = 57 else
"110111011111" when X = 70 AND Y = 57 else
"110111011111" when X = 71 AND Y = 57 else
"110111011111" when X = 72 AND Y = 57 else
"110111011111" when X = 73 AND Y = 57 else
"110111011111" when X = 74 AND Y = 57 else
"110111011111" when X = 75 AND Y = 57 else
"110111011111" when X = 76 AND Y = 57 else
"110111011111" when X = 77 AND Y = 57 else
"110111011111" when X = 78 AND Y = 57 else
"110111011111" when X = 79 AND Y = 57 else
"110111011111" when X = 80 AND Y = 57 else
"110111011111" when X = 81 AND Y = 57 else
"110111011111" when X = 82 AND Y = 57 else
"110111011111" when X = 83 AND Y = 57 else
"110111011111" when X = 84 AND Y = 57 else
"110111011111" when X = 85 AND Y = 57 else
"110111011111" when X = 86 AND Y = 57 else
"110111011111" when X = 87 AND Y = 57 else
"110111011111" when X = 88 AND Y = 57 else
"110111011111" when X = 89 AND Y = 57 else
"110111011111" when X = 90 AND Y = 57 else
"110111011111" when X = 91 AND Y = 57 else
"110111011111" when X = 92 AND Y = 57 else
"110111011111" when X = 93 AND Y = 57 else
"110111011111" when X = 94 AND Y = 57 else
"111111111111" when X = 95 AND Y = 57 else
"111111111111" when X = 96 AND Y = 57 else
"111111111111" when X = 97 AND Y = 57 else
"111111111111" when X = 98 AND Y = 57 else
"111111111111" when X = 99 AND Y = 57 else
"111111111111" when X = 100 AND Y = 57 else
"111111111111" when X = 101 AND Y = 57 else
"111111111111" when X = 102 AND Y = 57 else
"111111111111" when X = 103 AND Y = 57 else
"111111111111" when X = 104 AND Y = 57 else
"111111111111" when X = 105 AND Y = 57 else
"111111111111" when X = 106 AND Y = 57 else
"111111111111" when X = 107 AND Y = 57 else
"111111111111" when X = 108 AND Y = 57 else
"111111111111" when X = 109 AND Y = 57 else
"111111111111" when X = 110 AND Y = 57 else
"111111111111" when X = 111 AND Y = 57 else
"111111111111" when X = 112 AND Y = 57 else
"111111111111" when X = 113 AND Y = 57 else
"111111111111" when X = 114 AND Y = 57 else
"111111111111" when X = 115 AND Y = 57 else
"111111111111" when X = 116 AND Y = 57 else
"111111111111" when X = 117 AND Y = 57 else
"111111111111" when X = 118 AND Y = 57 else
"111111111111" when X = 119 AND Y = 57 else
"111111111111" when X = 120 AND Y = 57 else
"111111111111" when X = 121 AND Y = 57 else
"111111111111" when X = 122 AND Y = 57 else
"111111111111" when X = 123 AND Y = 57 else
"111111111111" when X = 124 AND Y = 57 else
"111111111111" when X = 125 AND Y = 57 else
"111111111111" when X = 126 AND Y = 57 else
"111111111111" when X = 127 AND Y = 57 else
"111111111111" when X = 128 AND Y = 57 else
"111111111111" when X = 129 AND Y = 57 else
"111111111111" when X = 130 AND Y = 57 else
"111111111111" when X = 131 AND Y = 57 else
"111111111111" when X = 132 AND Y = 57 else
"111111111111" when X = 133 AND Y = 57 else
"111111111111" when X = 134 AND Y = 57 else
"111111111111" when X = 135 AND Y = 57 else
"111111111111" when X = 136 AND Y = 57 else
"111111111111" when X = 137 AND Y = 57 else
"111111111111" when X = 138 AND Y = 57 else
"111111111111" when X = 139 AND Y = 57 else
"111111111111" when X = 140 AND Y = 57 else
"111111111111" when X = 141 AND Y = 57 else
"111111111111" when X = 142 AND Y = 57 else
"111111111111" when X = 143 AND Y = 57 else
"111111111111" when X = 144 AND Y = 57 else
"111111111111" when X = 145 AND Y = 57 else
"111111111111" when X = 146 AND Y = 57 else
"111111111111" when X = 147 AND Y = 57 else
"111111111111" when X = 148 AND Y = 57 else
"111111111111" when X = 149 AND Y = 57 else
"111111111111" when X = 150 AND Y = 57 else
"111111111111" when X = 151 AND Y = 57 else
"111111111111" when X = 152 AND Y = 57 else
"111111111111" when X = 153 AND Y = 57 else
"111111111111" when X = 154 AND Y = 57 else
"111111111111" when X = 155 AND Y = 57 else
"111111111111" when X = 156 AND Y = 57 else
"111111111111" when X = 157 AND Y = 57 else
"111111111111" when X = 158 AND Y = 57 else
"111111111111" when X = 159 AND Y = 57 else
"111111111111" when X = 160 AND Y = 57 else
"111111111111" when X = 161 AND Y = 57 else
"111111111111" when X = 162 AND Y = 57 else
"111111111111" when X = 163 AND Y = 57 else
"111111111111" when X = 164 AND Y = 57 else
"111111111111" when X = 165 AND Y = 57 else
"111111111111" when X = 166 AND Y = 57 else
"111111111111" when X = 167 AND Y = 57 else
"111111111111" when X = 168 AND Y = 57 else
"111111111111" when X = 169 AND Y = 57 else
"111111111111" when X = 170 AND Y = 57 else
"111111111111" when X = 171 AND Y = 57 else
"111111111111" when X = 172 AND Y = 57 else
"111111111111" when X = 173 AND Y = 57 else
"111111111111" when X = 174 AND Y = 57 else
"111111111111" when X = 175 AND Y = 57 else
"111111111111" when X = 176 AND Y = 57 else
"111111111111" when X = 177 AND Y = 57 else
"111111111111" when X = 178 AND Y = 57 else
"111111111111" when X = 179 AND Y = 57 else
"111111111111" when X = 180 AND Y = 57 else
"111111111111" when X = 181 AND Y = 57 else
"111111111111" when X = 182 AND Y = 57 else
"111111111111" when X = 183 AND Y = 57 else
"111111111111" when X = 184 AND Y = 57 else
"111111111111" when X = 185 AND Y = 57 else
"111111111111" when X = 186 AND Y = 57 else
"111111111111" when X = 187 AND Y = 57 else
"111111111111" when X = 188 AND Y = 57 else
"111111111111" when X = 189 AND Y = 57 else
"111111111111" when X = 190 AND Y = 57 else
"111111111111" when X = 191 AND Y = 57 else
"111111111111" when X = 192 AND Y = 57 else
"111111111111" when X = 193 AND Y = 57 else
"111111111111" when X = 194 AND Y = 57 else
"111111111111" when X = 195 AND Y = 57 else
"111111111111" when X = 196 AND Y = 57 else
"111111111111" when X = 197 AND Y = 57 else
"111111111111" when X = 198 AND Y = 57 else
"111111111111" when X = 199 AND Y = 57 else
"111111111111" when X = 200 AND Y = 57 else
"111111111111" when X = 201 AND Y = 57 else
"111111111111" when X = 202 AND Y = 57 else
"111111111111" when X = 203 AND Y = 57 else
"111111111111" when X = 204 AND Y = 57 else
"111111111111" when X = 205 AND Y = 57 else
"111111111111" when X = 206 AND Y = 57 else
"111111111111" when X = 207 AND Y = 57 else
"111111111111" when X = 208 AND Y = 57 else
"111111111111" when X = 209 AND Y = 57 else
"111111111111" when X = 210 AND Y = 57 else
"111111111111" when X = 211 AND Y = 57 else
"111111111111" when X = 212 AND Y = 57 else
"111111111111" when X = 213 AND Y = 57 else
"111111111111" when X = 214 AND Y = 57 else
"111111111111" when X = 215 AND Y = 57 else
"111111111111" when X = 216 AND Y = 57 else
"111111111111" when X = 217 AND Y = 57 else
"111111111111" when X = 218 AND Y = 57 else
"111111111111" when X = 219 AND Y = 57 else
"111111111111" when X = 220 AND Y = 57 else
"111111111111" when X = 221 AND Y = 57 else
"111111111111" when X = 222 AND Y = 57 else
"111111111111" when X = 223 AND Y = 57 else
"111111111111" when X = 224 AND Y = 57 else
"111111111111" when X = 225 AND Y = 57 else
"111111111111" when X = 226 AND Y = 57 else
"111111111111" when X = 227 AND Y = 57 else
"111111111111" when X = 228 AND Y = 57 else
"111111111111" when X = 229 AND Y = 57 else
"111111111111" when X = 230 AND Y = 57 else
"111111111111" when X = 231 AND Y = 57 else
"111111111111" when X = 232 AND Y = 57 else
"111111111111" when X = 233 AND Y = 57 else
"111111111111" when X = 234 AND Y = 57 else
"111111111111" when X = 235 AND Y = 57 else
"111111111111" when X = 236 AND Y = 57 else
"111111111111" when X = 237 AND Y = 57 else
"111111111111" when X = 238 AND Y = 57 else
"111111111111" when X = 239 AND Y = 57 else
"111111111111" when X = 240 AND Y = 57 else
"111111111111" when X = 241 AND Y = 57 else
"111111111111" when X = 242 AND Y = 57 else
"111111111111" when X = 243 AND Y = 57 else
"111111111111" when X = 244 AND Y = 57 else
"111111111111" when X = 245 AND Y = 57 else
"111111111111" when X = 246 AND Y = 57 else
"111111111111" when X = 247 AND Y = 57 else
"111111111111" when X = 248 AND Y = 57 else
"111111111111" when X = 249 AND Y = 57 else
"111111111111" when X = 250 AND Y = 57 else
"111111111111" when X = 251 AND Y = 57 else
"111111111111" when X = 252 AND Y = 57 else
"111111111111" when X = 253 AND Y = 57 else
"111111111111" when X = 254 AND Y = 57 else
"111111111111" when X = 255 AND Y = 57 else
"111111111111" when X = 256 AND Y = 57 else
"111111111111" when X = 257 AND Y = 57 else
"111111111111" when X = 258 AND Y = 57 else
"111111111111" when X = 259 AND Y = 57 else
"111111111111" when X = 260 AND Y = 57 else
"111111111111" when X = 261 AND Y = 57 else
"111111111111" when X = 262 AND Y = 57 else
"111111111111" when X = 263 AND Y = 57 else
"111111111111" when X = 264 AND Y = 57 else
"110111011111" when X = 265 AND Y = 57 else
"110111011111" when X = 266 AND Y = 57 else
"110111011111" when X = 267 AND Y = 57 else
"110111011111" when X = 268 AND Y = 57 else
"110111011111" when X = 269 AND Y = 57 else
"110111011111" when X = 270 AND Y = 57 else
"110111011111" when X = 271 AND Y = 57 else
"110111011111" when X = 272 AND Y = 57 else
"110111011111" when X = 273 AND Y = 57 else
"110111011111" when X = 274 AND Y = 57 else
"110111011111" when X = 275 AND Y = 57 else
"110111011111" when X = 276 AND Y = 57 else
"110111011111" when X = 277 AND Y = 57 else
"110111011111" when X = 278 AND Y = 57 else
"110111011111" when X = 279 AND Y = 57 else
"000000000000" when X = 280 AND Y = 57 else
"000000000000" when X = 281 AND Y = 57 else
"000000000000" when X = 282 AND Y = 57 else
"000000000000" when X = 283 AND Y = 57 else
"000000000000" when X = 284 AND Y = 57 else
"000000000000" when X = 285 AND Y = 57 else
"000000000000" when X = 286 AND Y = 57 else
"000000000000" when X = 287 AND Y = 57 else
"000000000000" when X = 288 AND Y = 57 else
"000000000000" when X = 289 AND Y = 57 else
"000000000000" when X = 290 AND Y = 57 else
"000000000000" when X = 291 AND Y = 57 else
"000000000000" when X = 292 AND Y = 57 else
"000000000000" when X = 293 AND Y = 57 else
"000000000000" when X = 294 AND Y = 57 else
"000000000000" when X = 295 AND Y = 57 else
"000000000000" when X = 296 AND Y = 57 else
"000000000000" when X = 297 AND Y = 57 else
"000000000000" when X = 298 AND Y = 57 else
"000000000000" when X = 299 AND Y = 57 else
"000000000000" when X = 300 AND Y = 57 else
"000000000000" when X = 301 AND Y = 57 else
"000000000000" when X = 302 AND Y = 57 else
"000000000000" when X = 303 AND Y = 57 else
"000000000000" when X = 304 AND Y = 57 else
"000000000000" when X = 305 AND Y = 57 else
"000000000000" when X = 306 AND Y = 57 else
"000000000000" when X = 307 AND Y = 57 else
"000000000000" when X = 308 AND Y = 57 else
"000000000000" when X = 309 AND Y = 57 else
"000000000000" when X = 310 AND Y = 57 else
"000000000000" when X = 311 AND Y = 57 else
"000000000000" when X = 312 AND Y = 57 else
"000000000000" when X = 313 AND Y = 57 else
"000000000000" when X = 314 AND Y = 57 else
"000000000000" when X = 315 AND Y = 57 else
"000000000000" when X = 316 AND Y = 57 else
"000000000000" when X = 317 AND Y = 57 else
"000000000000" when X = 318 AND Y = 57 else
"000000000000" when X = 319 AND Y = 57 else
"000000000000" when X = 320 AND Y = 57 else
"000000000000" when X = 321 AND Y = 57 else
"000000000000" when X = 322 AND Y = 57 else
"000000000000" when X = 323 AND Y = 57 else
"000000000000" when X = 324 AND Y = 57 else
"100010011101" when X = 0 AND Y = 58 else
"100010011101" when X = 1 AND Y = 58 else
"100010011101" when X = 2 AND Y = 58 else
"100010011101" when X = 3 AND Y = 58 else
"100010011101" when X = 4 AND Y = 58 else
"100010011101" when X = 5 AND Y = 58 else
"100010011101" when X = 6 AND Y = 58 else
"100010011101" when X = 7 AND Y = 58 else
"100010011101" when X = 8 AND Y = 58 else
"100010011101" when X = 9 AND Y = 58 else
"100010011101" when X = 10 AND Y = 58 else
"100010011101" when X = 11 AND Y = 58 else
"100010011101" when X = 12 AND Y = 58 else
"100010011101" when X = 13 AND Y = 58 else
"100010011101" when X = 14 AND Y = 58 else
"100010011101" when X = 15 AND Y = 58 else
"100010011101" when X = 16 AND Y = 58 else
"100010011101" when X = 17 AND Y = 58 else
"100010011101" when X = 18 AND Y = 58 else
"100010011101" when X = 19 AND Y = 58 else
"100010011101" when X = 20 AND Y = 58 else
"100010011101" when X = 21 AND Y = 58 else
"100010011101" when X = 22 AND Y = 58 else
"100010011101" when X = 23 AND Y = 58 else
"100010011101" when X = 24 AND Y = 58 else
"100010011101" when X = 25 AND Y = 58 else
"100010011101" when X = 26 AND Y = 58 else
"100010011101" when X = 27 AND Y = 58 else
"100010011101" when X = 28 AND Y = 58 else
"100010011101" when X = 29 AND Y = 58 else
"100010011101" when X = 30 AND Y = 58 else
"100010011101" when X = 31 AND Y = 58 else
"100010011101" when X = 32 AND Y = 58 else
"100010011101" when X = 33 AND Y = 58 else
"100010011101" when X = 34 AND Y = 58 else
"100010011101" when X = 35 AND Y = 58 else
"100010011101" when X = 36 AND Y = 58 else
"100010011101" when X = 37 AND Y = 58 else
"100010011101" when X = 38 AND Y = 58 else
"100010011101" when X = 39 AND Y = 58 else
"110111011111" when X = 40 AND Y = 58 else
"110111011111" when X = 41 AND Y = 58 else
"110111011111" when X = 42 AND Y = 58 else
"110111011111" when X = 43 AND Y = 58 else
"110111011111" when X = 44 AND Y = 58 else
"110111011111" when X = 45 AND Y = 58 else
"110111011111" when X = 46 AND Y = 58 else
"110111011111" when X = 47 AND Y = 58 else
"110111011111" when X = 48 AND Y = 58 else
"110111011111" when X = 49 AND Y = 58 else
"110111011111" when X = 50 AND Y = 58 else
"110111011111" when X = 51 AND Y = 58 else
"110111011111" when X = 52 AND Y = 58 else
"110111011111" when X = 53 AND Y = 58 else
"110111011111" when X = 54 AND Y = 58 else
"110111011111" when X = 55 AND Y = 58 else
"110111011111" when X = 56 AND Y = 58 else
"110111011111" when X = 57 AND Y = 58 else
"110111011111" when X = 58 AND Y = 58 else
"110111011111" when X = 59 AND Y = 58 else
"110111011111" when X = 60 AND Y = 58 else
"110111011111" when X = 61 AND Y = 58 else
"110111011111" when X = 62 AND Y = 58 else
"110111011111" when X = 63 AND Y = 58 else
"110111011111" when X = 64 AND Y = 58 else
"110111011111" when X = 65 AND Y = 58 else
"110111011111" when X = 66 AND Y = 58 else
"110111011111" when X = 67 AND Y = 58 else
"110111011111" when X = 68 AND Y = 58 else
"110111011111" when X = 69 AND Y = 58 else
"110111011111" when X = 70 AND Y = 58 else
"110111011111" when X = 71 AND Y = 58 else
"110111011111" when X = 72 AND Y = 58 else
"110111011111" when X = 73 AND Y = 58 else
"110111011111" when X = 74 AND Y = 58 else
"110111011111" when X = 75 AND Y = 58 else
"110111011111" when X = 76 AND Y = 58 else
"110111011111" when X = 77 AND Y = 58 else
"110111011111" when X = 78 AND Y = 58 else
"110111011111" when X = 79 AND Y = 58 else
"110111011111" when X = 80 AND Y = 58 else
"110111011111" when X = 81 AND Y = 58 else
"110111011111" when X = 82 AND Y = 58 else
"110111011111" when X = 83 AND Y = 58 else
"110111011111" when X = 84 AND Y = 58 else
"110111011111" when X = 85 AND Y = 58 else
"110111011111" when X = 86 AND Y = 58 else
"110111011111" when X = 87 AND Y = 58 else
"110111011111" when X = 88 AND Y = 58 else
"110111011111" when X = 89 AND Y = 58 else
"110111011111" when X = 90 AND Y = 58 else
"110111011111" when X = 91 AND Y = 58 else
"110111011111" when X = 92 AND Y = 58 else
"110111011111" when X = 93 AND Y = 58 else
"110111011111" when X = 94 AND Y = 58 else
"111111111111" when X = 95 AND Y = 58 else
"111111111111" when X = 96 AND Y = 58 else
"111111111111" when X = 97 AND Y = 58 else
"111111111111" when X = 98 AND Y = 58 else
"111111111111" when X = 99 AND Y = 58 else
"111111111111" when X = 100 AND Y = 58 else
"111111111111" when X = 101 AND Y = 58 else
"111111111111" when X = 102 AND Y = 58 else
"111111111111" when X = 103 AND Y = 58 else
"111111111111" when X = 104 AND Y = 58 else
"111111111111" when X = 105 AND Y = 58 else
"111111111111" when X = 106 AND Y = 58 else
"111111111111" when X = 107 AND Y = 58 else
"111111111111" when X = 108 AND Y = 58 else
"111111111111" when X = 109 AND Y = 58 else
"111111111111" when X = 110 AND Y = 58 else
"111111111111" when X = 111 AND Y = 58 else
"111111111111" when X = 112 AND Y = 58 else
"111111111111" when X = 113 AND Y = 58 else
"111111111111" when X = 114 AND Y = 58 else
"111111111111" when X = 115 AND Y = 58 else
"111111111111" when X = 116 AND Y = 58 else
"111111111111" when X = 117 AND Y = 58 else
"111111111111" when X = 118 AND Y = 58 else
"111111111111" when X = 119 AND Y = 58 else
"111111111111" when X = 120 AND Y = 58 else
"111111111111" when X = 121 AND Y = 58 else
"111111111111" when X = 122 AND Y = 58 else
"111111111111" when X = 123 AND Y = 58 else
"111111111111" when X = 124 AND Y = 58 else
"111111111111" when X = 125 AND Y = 58 else
"111111111111" when X = 126 AND Y = 58 else
"111111111111" when X = 127 AND Y = 58 else
"111111111111" when X = 128 AND Y = 58 else
"111111111111" when X = 129 AND Y = 58 else
"111111111111" when X = 130 AND Y = 58 else
"111111111111" when X = 131 AND Y = 58 else
"111111111111" when X = 132 AND Y = 58 else
"111111111111" when X = 133 AND Y = 58 else
"111111111111" when X = 134 AND Y = 58 else
"111111111111" when X = 135 AND Y = 58 else
"111111111111" when X = 136 AND Y = 58 else
"111111111111" when X = 137 AND Y = 58 else
"111111111111" when X = 138 AND Y = 58 else
"111111111111" when X = 139 AND Y = 58 else
"111111111111" when X = 140 AND Y = 58 else
"111111111111" when X = 141 AND Y = 58 else
"111111111111" when X = 142 AND Y = 58 else
"111111111111" when X = 143 AND Y = 58 else
"111111111111" when X = 144 AND Y = 58 else
"111111111111" when X = 145 AND Y = 58 else
"111111111111" when X = 146 AND Y = 58 else
"111111111111" when X = 147 AND Y = 58 else
"111111111111" when X = 148 AND Y = 58 else
"111111111111" when X = 149 AND Y = 58 else
"111111111111" when X = 150 AND Y = 58 else
"111111111111" when X = 151 AND Y = 58 else
"111111111111" when X = 152 AND Y = 58 else
"111111111111" when X = 153 AND Y = 58 else
"111111111111" when X = 154 AND Y = 58 else
"111111111111" when X = 155 AND Y = 58 else
"111111111111" when X = 156 AND Y = 58 else
"111111111111" when X = 157 AND Y = 58 else
"111111111111" when X = 158 AND Y = 58 else
"111111111111" when X = 159 AND Y = 58 else
"111111111111" when X = 160 AND Y = 58 else
"111111111111" when X = 161 AND Y = 58 else
"111111111111" when X = 162 AND Y = 58 else
"111111111111" when X = 163 AND Y = 58 else
"111111111111" when X = 164 AND Y = 58 else
"111111111111" when X = 165 AND Y = 58 else
"111111111111" when X = 166 AND Y = 58 else
"111111111111" when X = 167 AND Y = 58 else
"111111111111" when X = 168 AND Y = 58 else
"111111111111" when X = 169 AND Y = 58 else
"111111111111" when X = 170 AND Y = 58 else
"111111111111" when X = 171 AND Y = 58 else
"111111111111" when X = 172 AND Y = 58 else
"111111111111" when X = 173 AND Y = 58 else
"111111111111" when X = 174 AND Y = 58 else
"111111111111" when X = 175 AND Y = 58 else
"111111111111" when X = 176 AND Y = 58 else
"111111111111" when X = 177 AND Y = 58 else
"111111111111" when X = 178 AND Y = 58 else
"111111111111" when X = 179 AND Y = 58 else
"111111111111" when X = 180 AND Y = 58 else
"111111111111" when X = 181 AND Y = 58 else
"111111111111" when X = 182 AND Y = 58 else
"111111111111" when X = 183 AND Y = 58 else
"111111111111" when X = 184 AND Y = 58 else
"111111111111" when X = 185 AND Y = 58 else
"111111111111" when X = 186 AND Y = 58 else
"111111111111" when X = 187 AND Y = 58 else
"111111111111" when X = 188 AND Y = 58 else
"111111111111" when X = 189 AND Y = 58 else
"111111111111" when X = 190 AND Y = 58 else
"111111111111" when X = 191 AND Y = 58 else
"111111111111" when X = 192 AND Y = 58 else
"111111111111" when X = 193 AND Y = 58 else
"111111111111" when X = 194 AND Y = 58 else
"111111111111" when X = 195 AND Y = 58 else
"111111111111" when X = 196 AND Y = 58 else
"111111111111" when X = 197 AND Y = 58 else
"111111111111" when X = 198 AND Y = 58 else
"111111111111" when X = 199 AND Y = 58 else
"111111111111" when X = 200 AND Y = 58 else
"111111111111" when X = 201 AND Y = 58 else
"111111111111" when X = 202 AND Y = 58 else
"111111111111" when X = 203 AND Y = 58 else
"111111111111" when X = 204 AND Y = 58 else
"111111111111" when X = 205 AND Y = 58 else
"111111111111" when X = 206 AND Y = 58 else
"111111111111" when X = 207 AND Y = 58 else
"111111111111" when X = 208 AND Y = 58 else
"111111111111" when X = 209 AND Y = 58 else
"111111111111" when X = 210 AND Y = 58 else
"111111111111" when X = 211 AND Y = 58 else
"111111111111" when X = 212 AND Y = 58 else
"111111111111" when X = 213 AND Y = 58 else
"111111111111" when X = 214 AND Y = 58 else
"111111111111" when X = 215 AND Y = 58 else
"111111111111" when X = 216 AND Y = 58 else
"111111111111" when X = 217 AND Y = 58 else
"111111111111" when X = 218 AND Y = 58 else
"111111111111" when X = 219 AND Y = 58 else
"111111111111" when X = 220 AND Y = 58 else
"111111111111" when X = 221 AND Y = 58 else
"111111111111" when X = 222 AND Y = 58 else
"111111111111" when X = 223 AND Y = 58 else
"111111111111" when X = 224 AND Y = 58 else
"111111111111" when X = 225 AND Y = 58 else
"111111111111" when X = 226 AND Y = 58 else
"111111111111" when X = 227 AND Y = 58 else
"111111111111" when X = 228 AND Y = 58 else
"111111111111" when X = 229 AND Y = 58 else
"111111111111" when X = 230 AND Y = 58 else
"111111111111" when X = 231 AND Y = 58 else
"111111111111" when X = 232 AND Y = 58 else
"111111111111" when X = 233 AND Y = 58 else
"111111111111" when X = 234 AND Y = 58 else
"111111111111" when X = 235 AND Y = 58 else
"111111111111" when X = 236 AND Y = 58 else
"111111111111" when X = 237 AND Y = 58 else
"111111111111" when X = 238 AND Y = 58 else
"111111111111" when X = 239 AND Y = 58 else
"111111111111" when X = 240 AND Y = 58 else
"111111111111" when X = 241 AND Y = 58 else
"111111111111" when X = 242 AND Y = 58 else
"111111111111" when X = 243 AND Y = 58 else
"111111111111" when X = 244 AND Y = 58 else
"111111111111" when X = 245 AND Y = 58 else
"111111111111" when X = 246 AND Y = 58 else
"111111111111" when X = 247 AND Y = 58 else
"111111111111" when X = 248 AND Y = 58 else
"111111111111" when X = 249 AND Y = 58 else
"111111111111" when X = 250 AND Y = 58 else
"111111111111" when X = 251 AND Y = 58 else
"111111111111" when X = 252 AND Y = 58 else
"111111111111" when X = 253 AND Y = 58 else
"111111111111" when X = 254 AND Y = 58 else
"111111111111" when X = 255 AND Y = 58 else
"111111111111" when X = 256 AND Y = 58 else
"111111111111" when X = 257 AND Y = 58 else
"111111111111" when X = 258 AND Y = 58 else
"111111111111" when X = 259 AND Y = 58 else
"111111111111" when X = 260 AND Y = 58 else
"111111111111" when X = 261 AND Y = 58 else
"111111111111" when X = 262 AND Y = 58 else
"111111111111" when X = 263 AND Y = 58 else
"111111111111" when X = 264 AND Y = 58 else
"110111011111" when X = 265 AND Y = 58 else
"110111011111" when X = 266 AND Y = 58 else
"110111011111" when X = 267 AND Y = 58 else
"110111011111" when X = 268 AND Y = 58 else
"110111011111" when X = 269 AND Y = 58 else
"110111011111" when X = 270 AND Y = 58 else
"110111011111" when X = 271 AND Y = 58 else
"110111011111" when X = 272 AND Y = 58 else
"110111011111" when X = 273 AND Y = 58 else
"110111011111" when X = 274 AND Y = 58 else
"110111011111" when X = 275 AND Y = 58 else
"110111011111" when X = 276 AND Y = 58 else
"110111011111" when X = 277 AND Y = 58 else
"110111011111" when X = 278 AND Y = 58 else
"110111011111" when X = 279 AND Y = 58 else
"000000000000" when X = 280 AND Y = 58 else
"000000000000" when X = 281 AND Y = 58 else
"000000000000" when X = 282 AND Y = 58 else
"000000000000" when X = 283 AND Y = 58 else
"000000000000" when X = 284 AND Y = 58 else
"000000000000" when X = 285 AND Y = 58 else
"000000000000" when X = 286 AND Y = 58 else
"000000000000" when X = 287 AND Y = 58 else
"000000000000" when X = 288 AND Y = 58 else
"000000000000" when X = 289 AND Y = 58 else
"000000000000" when X = 290 AND Y = 58 else
"000000000000" when X = 291 AND Y = 58 else
"000000000000" when X = 292 AND Y = 58 else
"000000000000" when X = 293 AND Y = 58 else
"000000000000" when X = 294 AND Y = 58 else
"000000000000" when X = 295 AND Y = 58 else
"000000000000" when X = 296 AND Y = 58 else
"000000000000" when X = 297 AND Y = 58 else
"000000000000" when X = 298 AND Y = 58 else
"000000000000" when X = 299 AND Y = 58 else
"000000000000" when X = 300 AND Y = 58 else
"000000000000" when X = 301 AND Y = 58 else
"000000000000" when X = 302 AND Y = 58 else
"000000000000" when X = 303 AND Y = 58 else
"000000000000" when X = 304 AND Y = 58 else
"000000000000" when X = 305 AND Y = 58 else
"000000000000" when X = 306 AND Y = 58 else
"000000000000" when X = 307 AND Y = 58 else
"000000000000" when X = 308 AND Y = 58 else
"000000000000" when X = 309 AND Y = 58 else
"000000000000" when X = 310 AND Y = 58 else
"000000000000" when X = 311 AND Y = 58 else
"000000000000" when X = 312 AND Y = 58 else
"000000000000" when X = 313 AND Y = 58 else
"000000000000" when X = 314 AND Y = 58 else
"000000000000" when X = 315 AND Y = 58 else
"000000000000" when X = 316 AND Y = 58 else
"000000000000" when X = 317 AND Y = 58 else
"000000000000" when X = 318 AND Y = 58 else
"000000000000" when X = 319 AND Y = 58 else
"000000000000" when X = 320 AND Y = 58 else
"000000000000" when X = 321 AND Y = 58 else
"000000000000" when X = 322 AND Y = 58 else
"000000000000" when X = 323 AND Y = 58 else
"000000000000" when X = 324 AND Y = 58 else
"100010011101" when X = 0 AND Y = 59 else
"100010011101" when X = 1 AND Y = 59 else
"100010011101" when X = 2 AND Y = 59 else
"100010011101" when X = 3 AND Y = 59 else
"100010011101" when X = 4 AND Y = 59 else
"100010011101" when X = 5 AND Y = 59 else
"100010011101" when X = 6 AND Y = 59 else
"100010011101" when X = 7 AND Y = 59 else
"100010011101" when X = 8 AND Y = 59 else
"100010011101" when X = 9 AND Y = 59 else
"100010011101" when X = 10 AND Y = 59 else
"100010011101" when X = 11 AND Y = 59 else
"100010011101" when X = 12 AND Y = 59 else
"100010011101" when X = 13 AND Y = 59 else
"100010011101" when X = 14 AND Y = 59 else
"100010011101" when X = 15 AND Y = 59 else
"100010011101" when X = 16 AND Y = 59 else
"100010011101" when X = 17 AND Y = 59 else
"100010011101" when X = 18 AND Y = 59 else
"100010011101" when X = 19 AND Y = 59 else
"100010011101" when X = 20 AND Y = 59 else
"100010011101" when X = 21 AND Y = 59 else
"100010011101" when X = 22 AND Y = 59 else
"100010011101" when X = 23 AND Y = 59 else
"100010011101" when X = 24 AND Y = 59 else
"100010011101" when X = 25 AND Y = 59 else
"100010011101" when X = 26 AND Y = 59 else
"100010011101" when X = 27 AND Y = 59 else
"100010011101" when X = 28 AND Y = 59 else
"100010011101" when X = 29 AND Y = 59 else
"100010011101" when X = 30 AND Y = 59 else
"100010011101" when X = 31 AND Y = 59 else
"100010011101" when X = 32 AND Y = 59 else
"100010011101" when X = 33 AND Y = 59 else
"100010011101" when X = 34 AND Y = 59 else
"100010011101" when X = 35 AND Y = 59 else
"100010011101" when X = 36 AND Y = 59 else
"100010011101" when X = 37 AND Y = 59 else
"100010011101" when X = 38 AND Y = 59 else
"100010011101" when X = 39 AND Y = 59 else
"110111011111" when X = 40 AND Y = 59 else
"110111011111" when X = 41 AND Y = 59 else
"110111011111" when X = 42 AND Y = 59 else
"110111011111" when X = 43 AND Y = 59 else
"110111011111" when X = 44 AND Y = 59 else
"110111011111" when X = 45 AND Y = 59 else
"110111011111" when X = 46 AND Y = 59 else
"110111011111" when X = 47 AND Y = 59 else
"110111011111" when X = 48 AND Y = 59 else
"110111011111" when X = 49 AND Y = 59 else
"110111011111" when X = 50 AND Y = 59 else
"110111011111" when X = 51 AND Y = 59 else
"110111011111" when X = 52 AND Y = 59 else
"110111011111" when X = 53 AND Y = 59 else
"110111011111" when X = 54 AND Y = 59 else
"110111011111" when X = 55 AND Y = 59 else
"110111011111" when X = 56 AND Y = 59 else
"110111011111" when X = 57 AND Y = 59 else
"110111011111" when X = 58 AND Y = 59 else
"110111011111" when X = 59 AND Y = 59 else
"110111011111" when X = 60 AND Y = 59 else
"110111011111" when X = 61 AND Y = 59 else
"110111011111" when X = 62 AND Y = 59 else
"110111011111" when X = 63 AND Y = 59 else
"110111011111" when X = 64 AND Y = 59 else
"110111011111" when X = 65 AND Y = 59 else
"110111011111" when X = 66 AND Y = 59 else
"110111011111" when X = 67 AND Y = 59 else
"110111011111" when X = 68 AND Y = 59 else
"110111011111" when X = 69 AND Y = 59 else
"110111011111" when X = 70 AND Y = 59 else
"110111011111" when X = 71 AND Y = 59 else
"110111011111" when X = 72 AND Y = 59 else
"110111011111" when X = 73 AND Y = 59 else
"110111011111" when X = 74 AND Y = 59 else
"110111011111" when X = 75 AND Y = 59 else
"110111011111" when X = 76 AND Y = 59 else
"110111011111" when X = 77 AND Y = 59 else
"110111011111" when X = 78 AND Y = 59 else
"110111011111" when X = 79 AND Y = 59 else
"110111011111" when X = 80 AND Y = 59 else
"110111011111" when X = 81 AND Y = 59 else
"110111011111" when X = 82 AND Y = 59 else
"110111011111" when X = 83 AND Y = 59 else
"110111011111" when X = 84 AND Y = 59 else
"110111011111" when X = 85 AND Y = 59 else
"110111011111" when X = 86 AND Y = 59 else
"110111011111" when X = 87 AND Y = 59 else
"110111011111" when X = 88 AND Y = 59 else
"110111011111" when X = 89 AND Y = 59 else
"110111011111" when X = 90 AND Y = 59 else
"110111011111" when X = 91 AND Y = 59 else
"110111011111" when X = 92 AND Y = 59 else
"110111011111" when X = 93 AND Y = 59 else
"110111011111" when X = 94 AND Y = 59 else
"111111111111" when X = 95 AND Y = 59 else
"111111111111" when X = 96 AND Y = 59 else
"111111111111" when X = 97 AND Y = 59 else
"111111111111" when X = 98 AND Y = 59 else
"111111111111" when X = 99 AND Y = 59 else
"111111111111" when X = 100 AND Y = 59 else
"111111111111" when X = 101 AND Y = 59 else
"111111111111" when X = 102 AND Y = 59 else
"111111111111" when X = 103 AND Y = 59 else
"111111111111" when X = 104 AND Y = 59 else
"111111111111" when X = 105 AND Y = 59 else
"111111111111" when X = 106 AND Y = 59 else
"111111111111" when X = 107 AND Y = 59 else
"111111111111" when X = 108 AND Y = 59 else
"111111111111" when X = 109 AND Y = 59 else
"111111111111" when X = 110 AND Y = 59 else
"111111111111" when X = 111 AND Y = 59 else
"111111111111" when X = 112 AND Y = 59 else
"111111111111" when X = 113 AND Y = 59 else
"111111111111" when X = 114 AND Y = 59 else
"111111111111" when X = 115 AND Y = 59 else
"111111111111" when X = 116 AND Y = 59 else
"111111111111" when X = 117 AND Y = 59 else
"111111111111" when X = 118 AND Y = 59 else
"111111111111" when X = 119 AND Y = 59 else
"111111111111" when X = 120 AND Y = 59 else
"111111111111" when X = 121 AND Y = 59 else
"111111111111" when X = 122 AND Y = 59 else
"111111111111" when X = 123 AND Y = 59 else
"111111111111" when X = 124 AND Y = 59 else
"111111111111" when X = 125 AND Y = 59 else
"111111111111" when X = 126 AND Y = 59 else
"111111111111" when X = 127 AND Y = 59 else
"111111111111" when X = 128 AND Y = 59 else
"111111111111" when X = 129 AND Y = 59 else
"111111111111" when X = 130 AND Y = 59 else
"111111111111" when X = 131 AND Y = 59 else
"111111111111" when X = 132 AND Y = 59 else
"111111111111" when X = 133 AND Y = 59 else
"111111111111" when X = 134 AND Y = 59 else
"111111111111" when X = 135 AND Y = 59 else
"111111111111" when X = 136 AND Y = 59 else
"111111111111" when X = 137 AND Y = 59 else
"111111111111" when X = 138 AND Y = 59 else
"111111111111" when X = 139 AND Y = 59 else
"111111111111" when X = 140 AND Y = 59 else
"111111111111" when X = 141 AND Y = 59 else
"111111111111" when X = 142 AND Y = 59 else
"111111111111" when X = 143 AND Y = 59 else
"111111111111" when X = 144 AND Y = 59 else
"111111111111" when X = 145 AND Y = 59 else
"111111111111" when X = 146 AND Y = 59 else
"111111111111" when X = 147 AND Y = 59 else
"111111111111" when X = 148 AND Y = 59 else
"111111111111" when X = 149 AND Y = 59 else
"111111111111" when X = 150 AND Y = 59 else
"111111111111" when X = 151 AND Y = 59 else
"111111111111" when X = 152 AND Y = 59 else
"111111111111" when X = 153 AND Y = 59 else
"111111111111" when X = 154 AND Y = 59 else
"111111111111" when X = 155 AND Y = 59 else
"111111111111" when X = 156 AND Y = 59 else
"111111111111" when X = 157 AND Y = 59 else
"111111111111" when X = 158 AND Y = 59 else
"111111111111" when X = 159 AND Y = 59 else
"111111111111" when X = 160 AND Y = 59 else
"111111111111" when X = 161 AND Y = 59 else
"111111111111" when X = 162 AND Y = 59 else
"111111111111" when X = 163 AND Y = 59 else
"111111111111" when X = 164 AND Y = 59 else
"111111111111" when X = 165 AND Y = 59 else
"111111111111" when X = 166 AND Y = 59 else
"111111111111" when X = 167 AND Y = 59 else
"111111111111" when X = 168 AND Y = 59 else
"111111111111" when X = 169 AND Y = 59 else
"111111111111" when X = 170 AND Y = 59 else
"111111111111" when X = 171 AND Y = 59 else
"111111111111" when X = 172 AND Y = 59 else
"111111111111" when X = 173 AND Y = 59 else
"111111111111" when X = 174 AND Y = 59 else
"111111111111" when X = 175 AND Y = 59 else
"111111111111" when X = 176 AND Y = 59 else
"111111111111" when X = 177 AND Y = 59 else
"111111111111" when X = 178 AND Y = 59 else
"111111111111" when X = 179 AND Y = 59 else
"111111111111" when X = 180 AND Y = 59 else
"111111111111" when X = 181 AND Y = 59 else
"111111111111" when X = 182 AND Y = 59 else
"111111111111" when X = 183 AND Y = 59 else
"111111111111" when X = 184 AND Y = 59 else
"111111111111" when X = 185 AND Y = 59 else
"111111111111" when X = 186 AND Y = 59 else
"111111111111" when X = 187 AND Y = 59 else
"111111111111" when X = 188 AND Y = 59 else
"111111111111" when X = 189 AND Y = 59 else
"111111111111" when X = 190 AND Y = 59 else
"111111111111" when X = 191 AND Y = 59 else
"111111111111" when X = 192 AND Y = 59 else
"111111111111" when X = 193 AND Y = 59 else
"111111111111" when X = 194 AND Y = 59 else
"111111111111" when X = 195 AND Y = 59 else
"111111111111" when X = 196 AND Y = 59 else
"111111111111" when X = 197 AND Y = 59 else
"111111111111" when X = 198 AND Y = 59 else
"111111111111" when X = 199 AND Y = 59 else
"111111111111" when X = 200 AND Y = 59 else
"111111111111" when X = 201 AND Y = 59 else
"111111111111" when X = 202 AND Y = 59 else
"111111111111" when X = 203 AND Y = 59 else
"111111111111" when X = 204 AND Y = 59 else
"111111111111" when X = 205 AND Y = 59 else
"111111111111" when X = 206 AND Y = 59 else
"111111111111" when X = 207 AND Y = 59 else
"111111111111" when X = 208 AND Y = 59 else
"111111111111" when X = 209 AND Y = 59 else
"111111111111" when X = 210 AND Y = 59 else
"111111111111" when X = 211 AND Y = 59 else
"111111111111" when X = 212 AND Y = 59 else
"111111111111" when X = 213 AND Y = 59 else
"111111111111" when X = 214 AND Y = 59 else
"111111111111" when X = 215 AND Y = 59 else
"111111111111" when X = 216 AND Y = 59 else
"111111111111" when X = 217 AND Y = 59 else
"111111111111" when X = 218 AND Y = 59 else
"111111111111" when X = 219 AND Y = 59 else
"111111111111" when X = 220 AND Y = 59 else
"111111111111" when X = 221 AND Y = 59 else
"111111111111" when X = 222 AND Y = 59 else
"111111111111" when X = 223 AND Y = 59 else
"111111111111" when X = 224 AND Y = 59 else
"111111111111" when X = 225 AND Y = 59 else
"111111111111" when X = 226 AND Y = 59 else
"111111111111" when X = 227 AND Y = 59 else
"111111111111" when X = 228 AND Y = 59 else
"111111111111" when X = 229 AND Y = 59 else
"111111111111" when X = 230 AND Y = 59 else
"111111111111" when X = 231 AND Y = 59 else
"111111111111" when X = 232 AND Y = 59 else
"111111111111" when X = 233 AND Y = 59 else
"111111111111" when X = 234 AND Y = 59 else
"111111111111" when X = 235 AND Y = 59 else
"111111111111" when X = 236 AND Y = 59 else
"111111111111" when X = 237 AND Y = 59 else
"111111111111" when X = 238 AND Y = 59 else
"111111111111" when X = 239 AND Y = 59 else
"111111111111" when X = 240 AND Y = 59 else
"111111111111" when X = 241 AND Y = 59 else
"111111111111" when X = 242 AND Y = 59 else
"111111111111" when X = 243 AND Y = 59 else
"111111111111" when X = 244 AND Y = 59 else
"111111111111" when X = 245 AND Y = 59 else
"111111111111" when X = 246 AND Y = 59 else
"111111111111" when X = 247 AND Y = 59 else
"111111111111" when X = 248 AND Y = 59 else
"111111111111" when X = 249 AND Y = 59 else
"111111111111" when X = 250 AND Y = 59 else
"111111111111" when X = 251 AND Y = 59 else
"111111111111" when X = 252 AND Y = 59 else
"111111111111" when X = 253 AND Y = 59 else
"111111111111" when X = 254 AND Y = 59 else
"111111111111" when X = 255 AND Y = 59 else
"111111111111" when X = 256 AND Y = 59 else
"111111111111" when X = 257 AND Y = 59 else
"111111111111" when X = 258 AND Y = 59 else
"111111111111" when X = 259 AND Y = 59 else
"111111111111" when X = 260 AND Y = 59 else
"111111111111" when X = 261 AND Y = 59 else
"111111111111" when X = 262 AND Y = 59 else
"111111111111" when X = 263 AND Y = 59 else
"111111111111" when X = 264 AND Y = 59 else
"110111011111" when X = 265 AND Y = 59 else
"110111011111" when X = 266 AND Y = 59 else
"110111011111" when X = 267 AND Y = 59 else
"110111011111" when X = 268 AND Y = 59 else
"110111011111" when X = 269 AND Y = 59 else
"110111011111" when X = 270 AND Y = 59 else
"110111011111" when X = 271 AND Y = 59 else
"110111011111" when X = 272 AND Y = 59 else
"110111011111" when X = 273 AND Y = 59 else
"110111011111" when X = 274 AND Y = 59 else
"110111011111" when X = 275 AND Y = 59 else
"110111011111" when X = 276 AND Y = 59 else
"110111011111" when X = 277 AND Y = 59 else
"110111011111" when X = 278 AND Y = 59 else
"110111011111" when X = 279 AND Y = 59 else
"000000000000" when X = 280 AND Y = 59 else
"000000000000" when X = 281 AND Y = 59 else
"000000000000" when X = 282 AND Y = 59 else
"000000000000" when X = 283 AND Y = 59 else
"000000000000" when X = 284 AND Y = 59 else
"000000000000" when X = 285 AND Y = 59 else
"000000000000" when X = 286 AND Y = 59 else
"000000000000" when X = 287 AND Y = 59 else
"000000000000" when X = 288 AND Y = 59 else
"000000000000" when X = 289 AND Y = 59 else
"000000000000" when X = 290 AND Y = 59 else
"000000000000" when X = 291 AND Y = 59 else
"000000000000" when X = 292 AND Y = 59 else
"000000000000" when X = 293 AND Y = 59 else
"000000000000" when X = 294 AND Y = 59 else
"000000000000" when X = 295 AND Y = 59 else
"000000000000" when X = 296 AND Y = 59 else
"000000000000" when X = 297 AND Y = 59 else
"000000000000" when X = 298 AND Y = 59 else
"000000000000" when X = 299 AND Y = 59 else
"000000000000" when X = 300 AND Y = 59 else
"000000000000" when X = 301 AND Y = 59 else
"000000000000" when X = 302 AND Y = 59 else
"000000000000" when X = 303 AND Y = 59 else
"000000000000" when X = 304 AND Y = 59 else
"000000000000" when X = 305 AND Y = 59 else
"000000000000" when X = 306 AND Y = 59 else
"000000000000" when X = 307 AND Y = 59 else
"000000000000" when X = 308 AND Y = 59 else
"000000000000" when X = 309 AND Y = 59 else
"000000000000" when X = 310 AND Y = 59 else
"000000000000" when X = 311 AND Y = 59 else
"000000000000" when X = 312 AND Y = 59 else
"000000000000" when X = 313 AND Y = 59 else
"000000000000" when X = 314 AND Y = 59 else
"000000000000" when X = 315 AND Y = 59 else
"000000000000" when X = 316 AND Y = 59 else
"000000000000" when X = 317 AND Y = 59 else
"000000000000" when X = 318 AND Y = 59 else
"000000000000" when X = 319 AND Y = 59 else
"000000000000" when X = 320 AND Y = 59 else
"000000000000" when X = 321 AND Y = 59 else
"000000000000" when X = 322 AND Y = 59 else
"000000000000" when X = 323 AND Y = 59 else
"000000000000" when X = 324 AND Y = 59 else
"100010011101" when X = 0 AND Y = 60 else
"100010011101" when X = 1 AND Y = 60 else
"100010011101" when X = 2 AND Y = 60 else
"100010011101" when X = 3 AND Y = 60 else
"100010011101" when X = 4 AND Y = 60 else
"100010011101" when X = 5 AND Y = 60 else
"100010011101" when X = 6 AND Y = 60 else
"100010011101" when X = 7 AND Y = 60 else
"100010011101" when X = 8 AND Y = 60 else
"100010011101" when X = 9 AND Y = 60 else
"100010011101" when X = 10 AND Y = 60 else
"100010011101" when X = 11 AND Y = 60 else
"100010011101" when X = 12 AND Y = 60 else
"100010011101" when X = 13 AND Y = 60 else
"100010011101" when X = 14 AND Y = 60 else
"100010011101" when X = 15 AND Y = 60 else
"100010011101" when X = 16 AND Y = 60 else
"100010011101" when X = 17 AND Y = 60 else
"100010011101" when X = 18 AND Y = 60 else
"100010011101" when X = 19 AND Y = 60 else
"100010011101" when X = 20 AND Y = 60 else
"100010011101" when X = 21 AND Y = 60 else
"100010011101" when X = 22 AND Y = 60 else
"100010011101" when X = 23 AND Y = 60 else
"100010011101" when X = 24 AND Y = 60 else
"100010011101" when X = 25 AND Y = 60 else
"100010011101" when X = 26 AND Y = 60 else
"100010011101" when X = 27 AND Y = 60 else
"100010011101" when X = 28 AND Y = 60 else
"100010011101" when X = 29 AND Y = 60 else
"100010011101" when X = 30 AND Y = 60 else
"100010011101" when X = 31 AND Y = 60 else
"100010011101" when X = 32 AND Y = 60 else
"100010011101" when X = 33 AND Y = 60 else
"100010011101" when X = 34 AND Y = 60 else
"110111011111" when X = 35 AND Y = 60 else
"110111011111" when X = 36 AND Y = 60 else
"110111011111" when X = 37 AND Y = 60 else
"110111011111" when X = 38 AND Y = 60 else
"110111011111" when X = 39 AND Y = 60 else
"110111011111" when X = 40 AND Y = 60 else
"110111011111" when X = 41 AND Y = 60 else
"110111011111" when X = 42 AND Y = 60 else
"110111011111" when X = 43 AND Y = 60 else
"110111011111" when X = 44 AND Y = 60 else
"110111011111" when X = 45 AND Y = 60 else
"110111011111" when X = 46 AND Y = 60 else
"110111011111" when X = 47 AND Y = 60 else
"110111011111" when X = 48 AND Y = 60 else
"110111011111" when X = 49 AND Y = 60 else
"110111011111" when X = 50 AND Y = 60 else
"110111011111" when X = 51 AND Y = 60 else
"110111011111" when X = 52 AND Y = 60 else
"110111011111" when X = 53 AND Y = 60 else
"110111011111" when X = 54 AND Y = 60 else
"110111011111" when X = 55 AND Y = 60 else
"110111011111" when X = 56 AND Y = 60 else
"110111011111" when X = 57 AND Y = 60 else
"110111011111" when X = 58 AND Y = 60 else
"110111011111" when X = 59 AND Y = 60 else
"110111011111" when X = 60 AND Y = 60 else
"110111011111" when X = 61 AND Y = 60 else
"110111011111" when X = 62 AND Y = 60 else
"110111011111" when X = 63 AND Y = 60 else
"110111011111" when X = 64 AND Y = 60 else
"110111011111" when X = 65 AND Y = 60 else
"110111011111" when X = 66 AND Y = 60 else
"110111011111" when X = 67 AND Y = 60 else
"110111011111" when X = 68 AND Y = 60 else
"110111011111" when X = 69 AND Y = 60 else
"110111011111" when X = 70 AND Y = 60 else
"110111011111" when X = 71 AND Y = 60 else
"110111011111" when X = 72 AND Y = 60 else
"110111011111" when X = 73 AND Y = 60 else
"110111011111" when X = 74 AND Y = 60 else
"110111011111" when X = 75 AND Y = 60 else
"110111011111" when X = 76 AND Y = 60 else
"110111011111" when X = 77 AND Y = 60 else
"110111011111" when X = 78 AND Y = 60 else
"110111011111" when X = 79 AND Y = 60 else
"110111011111" when X = 80 AND Y = 60 else
"110111011111" when X = 81 AND Y = 60 else
"110111011111" when X = 82 AND Y = 60 else
"110111011111" when X = 83 AND Y = 60 else
"110111011111" when X = 84 AND Y = 60 else
"110111011111" when X = 85 AND Y = 60 else
"110111011111" when X = 86 AND Y = 60 else
"110111011111" when X = 87 AND Y = 60 else
"110111011111" when X = 88 AND Y = 60 else
"110111011111" when X = 89 AND Y = 60 else
"110111011111" when X = 90 AND Y = 60 else
"110111011111" when X = 91 AND Y = 60 else
"110111011111" when X = 92 AND Y = 60 else
"110111011111" when X = 93 AND Y = 60 else
"110111011111" when X = 94 AND Y = 60 else
"110111011111" when X = 95 AND Y = 60 else
"110111011111" when X = 96 AND Y = 60 else
"110111011111" when X = 97 AND Y = 60 else
"110111011111" when X = 98 AND Y = 60 else
"110111011111" when X = 99 AND Y = 60 else
"111111111111" when X = 100 AND Y = 60 else
"111111111111" when X = 101 AND Y = 60 else
"111111111111" when X = 102 AND Y = 60 else
"111111111111" when X = 103 AND Y = 60 else
"111111111111" when X = 104 AND Y = 60 else
"111111111111" when X = 105 AND Y = 60 else
"111111111111" when X = 106 AND Y = 60 else
"111111111111" when X = 107 AND Y = 60 else
"111111111111" when X = 108 AND Y = 60 else
"111111111111" when X = 109 AND Y = 60 else
"111111111111" when X = 110 AND Y = 60 else
"111111111111" when X = 111 AND Y = 60 else
"111111111111" when X = 112 AND Y = 60 else
"111111111111" when X = 113 AND Y = 60 else
"111111111111" when X = 114 AND Y = 60 else
"111111111111" when X = 115 AND Y = 60 else
"111111111111" when X = 116 AND Y = 60 else
"111111111111" when X = 117 AND Y = 60 else
"111111111111" when X = 118 AND Y = 60 else
"111111111111" when X = 119 AND Y = 60 else
"111111111111" when X = 120 AND Y = 60 else
"111111111111" when X = 121 AND Y = 60 else
"111111111111" when X = 122 AND Y = 60 else
"111111111111" when X = 123 AND Y = 60 else
"111111111111" when X = 124 AND Y = 60 else
"111111111111" when X = 125 AND Y = 60 else
"111111111111" when X = 126 AND Y = 60 else
"111111111111" when X = 127 AND Y = 60 else
"111111111111" when X = 128 AND Y = 60 else
"111111111111" when X = 129 AND Y = 60 else
"111111111111" when X = 130 AND Y = 60 else
"111111111111" when X = 131 AND Y = 60 else
"111111111111" when X = 132 AND Y = 60 else
"111111111111" when X = 133 AND Y = 60 else
"111111111111" when X = 134 AND Y = 60 else
"111111111111" when X = 135 AND Y = 60 else
"111111111111" when X = 136 AND Y = 60 else
"111111111111" when X = 137 AND Y = 60 else
"111111111111" when X = 138 AND Y = 60 else
"111111111111" when X = 139 AND Y = 60 else
"111111111111" when X = 140 AND Y = 60 else
"111111111111" when X = 141 AND Y = 60 else
"111111111111" when X = 142 AND Y = 60 else
"111111111111" when X = 143 AND Y = 60 else
"111111111111" when X = 144 AND Y = 60 else
"111111111111" when X = 145 AND Y = 60 else
"111111111111" when X = 146 AND Y = 60 else
"111111111111" when X = 147 AND Y = 60 else
"111111111111" when X = 148 AND Y = 60 else
"111111111111" when X = 149 AND Y = 60 else
"111111111111" when X = 150 AND Y = 60 else
"111111111111" when X = 151 AND Y = 60 else
"111111111111" when X = 152 AND Y = 60 else
"111111111111" when X = 153 AND Y = 60 else
"111111111111" when X = 154 AND Y = 60 else
"111111111111" when X = 155 AND Y = 60 else
"111111111111" when X = 156 AND Y = 60 else
"111111111111" when X = 157 AND Y = 60 else
"111111111111" when X = 158 AND Y = 60 else
"111111111111" when X = 159 AND Y = 60 else
"111111111111" when X = 160 AND Y = 60 else
"111111111111" when X = 161 AND Y = 60 else
"111111111111" when X = 162 AND Y = 60 else
"111111111111" when X = 163 AND Y = 60 else
"111111111111" when X = 164 AND Y = 60 else
"111111111111" when X = 165 AND Y = 60 else
"111111111111" when X = 166 AND Y = 60 else
"111111111111" when X = 167 AND Y = 60 else
"111111111111" when X = 168 AND Y = 60 else
"111111111111" when X = 169 AND Y = 60 else
"111111111111" when X = 170 AND Y = 60 else
"111111111111" when X = 171 AND Y = 60 else
"111111111111" when X = 172 AND Y = 60 else
"111111111111" when X = 173 AND Y = 60 else
"111111111111" when X = 174 AND Y = 60 else
"111111111111" when X = 175 AND Y = 60 else
"111111111111" when X = 176 AND Y = 60 else
"111111111111" when X = 177 AND Y = 60 else
"111111111111" when X = 178 AND Y = 60 else
"111111111111" when X = 179 AND Y = 60 else
"111111111111" when X = 180 AND Y = 60 else
"111111111111" when X = 181 AND Y = 60 else
"111111111111" when X = 182 AND Y = 60 else
"111111111111" when X = 183 AND Y = 60 else
"111111111111" when X = 184 AND Y = 60 else
"111111111111" when X = 185 AND Y = 60 else
"111111111111" when X = 186 AND Y = 60 else
"111111111111" when X = 187 AND Y = 60 else
"111111111111" when X = 188 AND Y = 60 else
"111111111111" when X = 189 AND Y = 60 else
"111111111111" when X = 190 AND Y = 60 else
"111111111111" when X = 191 AND Y = 60 else
"111111111111" when X = 192 AND Y = 60 else
"111111111111" when X = 193 AND Y = 60 else
"111111111111" when X = 194 AND Y = 60 else
"111111111111" when X = 195 AND Y = 60 else
"111111111111" when X = 196 AND Y = 60 else
"111111111111" when X = 197 AND Y = 60 else
"111111111111" when X = 198 AND Y = 60 else
"111111111111" when X = 199 AND Y = 60 else
"111111111111" when X = 200 AND Y = 60 else
"111111111111" when X = 201 AND Y = 60 else
"111111111111" when X = 202 AND Y = 60 else
"111111111111" when X = 203 AND Y = 60 else
"111111111111" when X = 204 AND Y = 60 else
"111111111111" when X = 205 AND Y = 60 else
"111111111111" when X = 206 AND Y = 60 else
"111111111111" when X = 207 AND Y = 60 else
"111111111111" when X = 208 AND Y = 60 else
"111111111111" when X = 209 AND Y = 60 else
"111111111111" when X = 210 AND Y = 60 else
"111111111111" when X = 211 AND Y = 60 else
"111111111111" when X = 212 AND Y = 60 else
"111111111111" when X = 213 AND Y = 60 else
"111111111111" when X = 214 AND Y = 60 else
"111111111111" when X = 215 AND Y = 60 else
"111111111111" when X = 216 AND Y = 60 else
"111111111111" when X = 217 AND Y = 60 else
"111111111111" when X = 218 AND Y = 60 else
"111111111111" when X = 219 AND Y = 60 else
"111111111111" when X = 220 AND Y = 60 else
"111111111111" when X = 221 AND Y = 60 else
"111111111111" when X = 222 AND Y = 60 else
"111111111111" when X = 223 AND Y = 60 else
"111111111111" when X = 224 AND Y = 60 else
"111111111111" when X = 225 AND Y = 60 else
"111111111111" when X = 226 AND Y = 60 else
"111111111111" when X = 227 AND Y = 60 else
"111111111111" when X = 228 AND Y = 60 else
"111111111111" when X = 229 AND Y = 60 else
"111111111111" when X = 230 AND Y = 60 else
"111111111111" when X = 231 AND Y = 60 else
"111111111111" when X = 232 AND Y = 60 else
"111111111111" when X = 233 AND Y = 60 else
"111111111111" when X = 234 AND Y = 60 else
"111111111111" when X = 235 AND Y = 60 else
"111111111111" when X = 236 AND Y = 60 else
"111111111111" when X = 237 AND Y = 60 else
"111111111111" when X = 238 AND Y = 60 else
"111111111111" when X = 239 AND Y = 60 else
"111111111111" when X = 240 AND Y = 60 else
"111111111111" when X = 241 AND Y = 60 else
"111111111111" when X = 242 AND Y = 60 else
"111111111111" when X = 243 AND Y = 60 else
"111111111111" when X = 244 AND Y = 60 else
"111111111111" when X = 245 AND Y = 60 else
"111111111111" when X = 246 AND Y = 60 else
"111111111111" when X = 247 AND Y = 60 else
"111111111111" when X = 248 AND Y = 60 else
"111111111111" when X = 249 AND Y = 60 else
"111111111111" when X = 250 AND Y = 60 else
"111111111111" when X = 251 AND Y = 60 else
"111111111111" when X = 252 AND Y = 60 else
"111111111111" when X = 253 AND Y = 60 else
"111111111111" when X = 254 AND Y = 60 else
"111111111111" when X = 255 AND Y = 60 else
"111111111111" when X = 256 AND Y = 60 else
"111111111111" when X = 257 AND Y = 60 else
"111111111111" when X = 258 AND Y = 60 else
"111111111111" when X = 259 AND Y = 60 else
"111111111111" when X = 260 AND Y = 60 else
"111111111111" when X = 261 AND Y = 60 else
"111111111111" when X = 262 AND Y = 60 else
"111111111111" when X = 263 AND Y = 60 else
"111111111111" when X = 264 AND Y = 60 else
"110111011111" when X = 265 AND Y = 60 else
"110111011111" when X = 266 AND Y = 60 else
"110111011111" when X = 267 AND Y = 60 else
"110111011111" when X = 268 AND Y = 60 else
"110111011111" when X = 269 AND Y = 60 else
"110111011111" when X = 270 AND Y = 60 else
"110111011111" when X = 271 AND Y = 60 else
"110111011111" when X = 272 AND Y = 60 else
"110111011111" when X = 273 AND Y = 60 else
"110111011111" when X = 274 AND Y = 60 else
"110111011111" when X = 275 AND Y = 60 else
"110111011111" when X = 276 AND Y = 60 else
"110111011111" when X = 277 AND Y = 60 else
"110111011111" when X = 278 AND Y = 60 else
"110111011111" when X = 279 AND Y = 60 else
"000000000000" when X = 280 AND Y = 60 else
"000000000000" when X = 281 AND Y = 60 else
"000000000000" when X = 282 AND Y = 60 else
"000000000000" when X = 283 AND Y = 60 else
"000000000000" when X = 284 AND Y = 60 else
"000000000000" when X = 285 AND Y = 60 else
"000000000000" when X = 286 AND Y = 60 else
"000000000000" when X = 287 AND Y = 60 else
"000000000000" when X = 288 AND Y = 60 else
"000000000000" when X = 289 AND Y = 60 else
"000000000000" when X = 290 AND Y = 60 else
"000000000000" when X = 291 AND Y = 60 else
"000000000000" when X = 292 AND Y = 60 else
"000000000000" when X = 293 AND Y = 60 else
"000000000000" when X = 294 AND Y = 60 else
"000000000000" when X = 295 AND Y = 60 else
"000000000000" when X = 296 AND Y = 60 else
"000000000000" when X = 297 AND Y = 60 else
"000000000000" when X = 298 AND Y = 60 else
"000000000000" when X = 299 AND Y = 60 else
"000000000000" when X = 300 AND Y = 60 else
"000000000000" when X = 301 AND Y = 60 else
"000000000000" when X = 302 AND Y = 60 else
"000000000000" when X = 303 AND Y = 60 else
"000000000000" when X = 304 AND Y = 60 else
"000000000000" when X = 305 AND Y = 60 else
"000000000000" when X = 306 AND Y = 60 else
"000000000000" when X = 307 AND Y = 60 else
"000000000000" when X = 308 AND Y = 60 else
"000000000000" when X = 309 AND Y = 60 else
"000000000000" when X = 310 AND Y = 60 else
"000000000000" when X = 311 AND Y = 60 else
"000000000000" when X = 312 AND Y = 60 else
"000000000000" when X = 313 AND Y = 60 else
"000000000000" when X = 314 AND Y = 60 else
"000000000000" when X = 315 AND Y = 60 else
"000000000000" when X = 316 AND Y = 60 else
"000000000000" when X = 317 AND Y = 60 else
"000000000000" when X = 318 AND Y = 60 else
"000000000000" when X = 319 AND Y = 60 else
"000000000000" when X = 320 AND Y = 60 else
"000000000000" when X = 321 AND Y = 60 else
"000000000000" when X = 322 AND Y = 60 else
"000000000000" when X = 323 AND Y = 60 else
"000000000000" when X = 324 AND Y = 60 else
"100010011101" when X = 0 AND Y = 61 else
"100010011101" when X = 1 AND Y = 61 else
"100010011101" when X = 2 AND Y = 61 else
"100010011101" when X = 3 AND Y = 61 else
"100010011101" when X = 4 AND Y = 61 else
"100010011101" when X = 5 AND Y = 61 else
"100010011101" when X = 6 AND Y = 61 else
"100010011101" when X = 7 AND Y = 61 else
"100010011101" when X = 8 AND Y = 61 else
"100010011101" when X = 9 AND Y = 61 else
"100010011101" when X = 10 AND Y = 61 else
"100010011101" when X = 11 AND Y = 61 else
"100010011101" when X = 12 AND Y = 61 else
"100010011101" when X = 13 AND Y = 61 else
"100010011101" when X = 14 AND Y = 61 else
"100010011101" when X = 15 AND Y = 61 else
"100010011101" when X = 16 AND Y = 61 else
"100010011101" when X = 17 AND Y = 61 else
"100010011101" when X = 18 AND Y = 61 else
"100010011101" when X = 19 AND Y = 61 else
"100010011101" when X = 20 AND Y = 61 else
"100010011101" when X = 21 AND Y = 61 else
"100010011101" when X = 22 AND Y = 61 else
"100010011101" when X = 23 AND Y = 61 else
"100010011101" when X = 24 AND Y = 61 else
"100010011101" when X = 25 AND Y = 61 else
"100010011101" when X = 26 AND Y = 61 else
"100010011101" when X = 27 AND Y = 61 else
"100010011101" when X = 28 AND Y = 61 else
"100010011101" when X = 29 AND Y = 61 else
"100010011101" when X = 30 AND Y = 61 else
"100010011101" when X = 31 AND Y = 61 else
"100010011101" when X = 32 AND Y = 61 else
"100010011101" when X = 33 AND Y = 61 else
"100010011101" when X = 34 AND Y = 61 else
"110111011111" when X = 35 AND Y = 61 else
"110111011111" when X = 36 AND Y = 61 else
"110111011111" when X = 37 AND Y = 61 else
"110111011111" when X = 38 AND Y = 61 else
"110111011111" when X = 39 AND Y = 61 else
"110111011111" when X = 40 AND Y = 61 else
"110111011111" when X = 41 AND Y = 61 else
"110111011111" when X = 42 AND Y = 61 else
"110111011111" when X = 43 AND Y = 61 else
"110111011111" when X = 44 AND Y = 61 else
"110111011111" when X = 45 AND Y = 61 else
"110111011111" when X = 46 AND Y = 61 else
"110111011111" when X = 47 AND Y = 61 else
"110111011111" when X = 48 AND Y = 61 else
"110111011111" when X = 49 AND Y = 61 else
"110111011111" when X = 50 AND Y = 61 else
"110111011111" when X = 51 AND Y = 61 else
"110111011111" when X = 52 AND Y = 61 else
"110111011111" when X = 53 AND Y = 61 else
"110111011111" when X = 54 AND Y = 61 else
"110111011111" when X = 55 AND Y = 61 else
"110111011111" when X = 56 AND Y = 61 else
"110111011111" when X = 57 AND Y = 61 else
"110111011111" when X = 58 AND Y = 61 else
"110111011111" when X = 59 AND Y = 61 else
"110111011111" when X = 60 AND Y = 61 else
"110111011111" when X = 61 AND Y = 61 else
"110111011111" when X = 62 AND Y = 61 else
"110111011111" when X = 63 AND Y = 61 else
"110111011111" when X = 64 AND Y = 61 else
"110111011111" when X = 65 AND Y = 61 else
"110111011111" when X = 66 AND Y = 61 else
"110111011111" when X = 67 AND Y = 61 else
"110111011111" when X = 68 AND Y = 61 else
"110111011111" when X = 69 AND Y = 61 else
"110111011111" when X = 70 AND Y = 61 else
"110111011111" when X = 71 AND Y = 61 else
"110111011111" when X = 72 AND Y = 61 else
"110111011111" when X = 73 AND Y = 61 else
"110111011111" when X = 74 AND Y = 61 else
"110111011111" when X = 75 AND Y = 61 else
"110111011111" when X = 76 AND Y = 61 else
"110111011111" when X = 77 AND Y = 61 else
"110111011111" when X = 78 AND Y = 61 else
"110111011111" when X = 79 AND Y = 61 else
"110111011111" when X = 80 AND Y = 61 else
"110111011111" when X = 81 AND Y = 61 else
"110111011111" when X = 82 AND Y = 61 else
"110111011111" when X = 83 AND Y = 61 else
"110111011111" when X = 84 AND Y = 61 else
"110111011111" when X = 85 AND Y = 61 else
"110111011111" when X = 86 AND Y = 61 else
"110111011111" when X = 87 AND Y = 61 else
"110111011111" when X = 88 AND Y = 61 else
"110111011111" when X = 89 AND Y = 61 else
"110111011111" when X = 90 AND Y = 61 else
"110111011111" when X = 91 AND Y = 61 else
"110111011111" when X = 92 AND Y = 61 else
"110111011111" when X = 93 AND Y = 61 else
"110111011111" when X = 94 AND Y = 61 else
"110111011111" when X = 95 AND Y = 61 else
"110111011111" when X = 96 AND Y = 61 else
"110111011111" when X = 97 AND Y = 61 else
"110111011111" when X = 98 AND Y = 61 else
"110111011111" when X = 99 AND Y = 61 else
"111111111111" when X = 100 AND Y = 61 else
"111111111111" when X = 101 AND Y = 61 else
"111111111111" when X = 102 AND Y = 61 else
"111111111111" when X = 103 AND Y = 61 else
"111111111111" when X = 104 AND Y = 61 else
"111111111111" when X = 105 AND Y = 61 else
"111111111111" when X = 106 AND Y = 61 else
"111111111111" when X = 107 AND Y = 61 else
"111111111111" when X = 108 AND Y = 61 else
"111111111111" when X = 109 AND Y = 61 else
"111111111111" when X = 110 AND Y = 61 else
"111111111111" when X = 111 AND Y = 61 else
"111111111111" when X = 112 AND Y = 61 else
"111111111111" when X = 113 AND Y = 61 else
"111111111111" when X = 114 AND Y = 61 else
"111111111111" when X = 115 AND Y = 61 else
"111111111111" when X = 116 AND Y = 61 else
"111111111111" when X = 117 AND Y = 61 else
"111111111111" when X = 118 AND Y = 61 else
"111111111111" when X = 119 AND Y = 61 else
"111111111111" when X = 120 AND Y = 61 else
"111111111111" when X = 121 AND Y = 61 else
"111111111111" when X = 122 AND Y = 61 else
"111111111111" when X = 123 AND Y = 61 else
"111111111111" when X = 124 AND Y = 61 else
"111111111111" when X = 125 AND Y = 61 else
"111111111111" when X = 126 AND Y = 61 else
"111111111111" when X = 127 AND Y = 61 else
"111111111111" when X = 128 AND Y = 61 else
"111111111111" when X = 129 AND Y = 61 else
"111111111111" when X = 130 AND Y = 61 else
"111111111111" when X = 131 AND Y = 61 else
"111111111111" when X = 132 AND Y = 61 else
"111111111111" when X = 133 AND Y = 61 else
"111111111111" when X = 134 AND Y = 61 else
"111111111111" when X = 135 AND Y = 61 else
"111111111111" when X = 136 AND Y = 61 else
"111111111111" when X = 137 AND Y = 61 else
"111111111111" when X = 138 AND Y = 61 else
"111111111111" when X = 139 AND Y = 61 else
"111111111111" when X = 140 AND Y = 61 else
"111111111111" when X = 141 AND Y = 61 else
"111111111111" when X = 142 AND Y = 61 else
"111111111111" when X = 143 AND Y = 61 else
"111111111111" when X = 144 AND Y = 61 else
"111111111111" when X = 145 AND Y = 61 else
"111111111111" when X = 146 AND Y = 61 else
"111111111111" when X = 147 AND Y = 61 else
"111111111111" when X = 148 AND Y = 61 else
"111111111111" when X = 149 AND Y = 61 else
"111111111111" when X = 150 AND Y = 61 else
"111111111111" when X = 151 AND Y = 61 else
"111111111111" when X = 152 AND Y = 61 else
"111111111111" when X = 153 AND Y = 61 else
"111111111111" when X = 154 AND Y = 61 else
"111111111111" when X = 155 AND Y = 61 else
"111111111111" when X = 156 AND Y = 61 else
"111111111111" when X = 157 AND Y = 61 else
"111111111111" when X = 158 AND Y = 61 else
"111111111111" when X = 159 AND Y = 61 else
"111111111111" when X = 160 AND Y = 61 else
"111111111111" when X = 161 AND Y = 61 else
"111111111111" when X = 162 AND Y = 61 else
"111111111111" when X = 163 AND Y = 61 else
"111111111111" when X = 164 AND Y = 61 else
"111111111111" when X = 165 AND Y = 61 else
"111111111111" when X = 166 AND Y = 61 else
"111111111111" when X = 167 AND Y = 61 else
"111111111111" when X = 168 AND Y = 61 else
"111111111111" when X = 169 AND Y = 61 else
"111111111111" when X = 170 AND Y = 61 else
"111111111111" when X = 171 AND Y = 61 else
"111111111111" when X = 172 AND Y = 61 else
"111111111111" when X = 173 AND Y = 61 else
"111111111111" when X = 174 AND Y = 61 else
"111111111111" when X = 175 AND Y = 61 else
"111111111111" when X = 176 AND Y = 61 else
"111111111111" when X = 177 AND Y = 61 else
"111111111111" when X = 178 AND Y = 61 else
"111111111111" when X = 179 AND Y = 61 else
"111111111111" when X = 180 AND Y = 61 else
"111111111111" when X = 181 AND Y = 61 else
"111111111111" when X = 182 AND Y = 61 else
"111111111111" when X = 183 AND Y = 61 else
"111111111111" when X = 184 AND Y = 61 else
"111111111111" when X = 185 AND Y = 61 else
"111111111111" when X = 186 AND Y = 61 else
"111111111111" when X = 187 AND Y = 61 else
"111111111111" when X = 188 AND Y = 61 else
"111111111111" when X = 189 AND Y = 61 else
"111111111111" when X = 190 AND Y = 61 else
"111111111111" when X = 191 AND Y = 61 else
"111111111111" when X = 192 AND Y = 61 else
"111111111111" when X = 193 AND Y = 61 else
"111111111111" when X = 194 AND Y = 61 else
"111111111111" when X = 195 AND Y = 61 else
"111111111111" when X = 196 AND Y = 61 else
"111111111111" when X = 197 AND Y = 61 else
"111111111111" when X = 198 AND Y = 61 else
"111111111111" when X = 199 AND Y = 61 else
"111111111111" when X = 200 AND Y = 61 else
"111111111111" when X = 201 AND Y = 61 else
"111111111111" when X = 202 AND Y = 61 else
"111111111111" when X = 203 AND Y = 61 else
"111111111111" when X = 204 AND Y = 61 else
"111111111111" when X = 205 AND Y = 61 else
"111111111111" when X = 206 AND Y = 61 else
"111111111111" when X = 207 AND Y = 61 else
"111111111111" when X = 208 AND Y = 61 else
"111111111111" when X = 209 AND Y = 61 else
"111111111111" when X = 210 AND Y = 61 else
"111111111111" when X = 211 AND Y = 61 else
"111111111111" when X = 212 AND Y = 61 else
"111111111111" when X = 213 AND Y = 61 else
"111111111111" when X = 214 AND Y = 61 else
"111111111111" when X = 215 AND Y = 61 else
"111111111111" when X = 216 AND Y = 61 else
"111111111111" when X = 217 AND Y = 61 else
"111111111111" when X = 218 AND Y = 61 else
"111111111111" when X = 219 AND Y = 61 else
"111111111111" when X = 220 AND Y = 61 else
"111111111111" when X = 221 AND Y = 61 else
"111111111111" when X = 222 AND Y = 61 else
"111111111111" when X = 223 AND Y = 61 else
"111111111111" when X = 224 AND Y = 61 else
"111111111111" when X = 225 AND Y = 61 else
"111111111111" when X = 226 AND Y = 61 else
"111111111111" when X = 227 AND Y = 61 else
"111111111111" when X = 228 AND Y = 61 else
"111111111111" when X = 229 AND Y = 61 else
"111111111111" when X = 230 AND Y = 61 else
"111111111111" when X = 231 AND Y = 61 else
"111111111111" when X = 232 AND Y = 61 else
"111111111111" when X = 233 AND Y = 61 else
"111111111111" when X = 234 AND Y = 61 else
"111111111111" when X = 235 AND Y = 61 else
"111111111111" when X = 236 AND Y = 61 else
"111111111111" when X = 237 AND Y = 61 else
"111111111111" when X = 238 AND Y = 61 else
"111111111111" when X = 239 AND Y = 61 else
"111111111111" when X = 240 AND Y = 61 else
"111111111111" when X = 241 AND Y = 61 else
"111111111111" when X = 242 AND Y = 61 else
"111111111111" when X = 243 AND Y = 61 else
"111111111111" when X = 244 AND Y = 61 else
"111111111111" when X = 245 AND Y = 61 else
"111111111111" when X = 246 AND Y = 61 else
"111111111111" when X = 247 AND Y = 61 else
"111111111111" when X = 248 AND Y = 61 else
"111111111111" when X = 249 AND Y = 61 else
"111111111111" when X = 250 AND Y = 61 else
"111111111111" when X = 251 AND Y = 61 else
"111111111111" when X = 252 AND Y = 61 else
"111111111111" when X = 253 AND Y = 61 else
"111111111111" when X = 254 AND Y = 61 else
"111111111111" when X = 255 AND Y = 61 else
"111111111111" when X = 256 AND Y = 61 else
"111111111111" when X = 257 AND Y = 61 else
"111111111111" when X = 258 AND Y = 61 else
"111111111111" when X = 259 AND Y = 61 else
"111111111111" when X = 260 AND Y = 61 else
"111111111111" when X = 261 AND Y = 61 else
"111111111111" when X = 262 AND Y = 61 else
"111111111111" when X = 263 AND Y = 61 else
"111111111111" when X = 264 AND Y = 61 else
"110111011111" when X = 265 AND Y = 61 else
"110111011111" when X = 266 AND Y = 61 else
"110111011111" when X = 267 AND Y = 61 else
"110111011111" when X = 268 AND Y = 61 else
"110111011111" when X = 269 AND Y = 61 else
"110111011111" when X = 270 AND Y = 61 else
"110111011111" when X = 271 AND Y = 61 else
"110111011111" when X = 272 AND Y = 61 else
"110111011111" when X = 273 AND Y = 61 else
"110111011111" when X = 274 AND Y = 61 else
"110111011111" when X = 275 AND Y = 61 else
"110111011111" when X = 276 AND Y = 61 else
"110111011111" when X = 277 AND Y = 61 else
"110111011111" when X = 278 AND Y = 61 else
"110111011111" when X = 279 AND Y = 61 else
"000000000000" when X = 280 AND Y = 61 else
"000000000000" when X = 281 AND Y = 61 else
"000000000000" when X = 282 AND Y = 61 else
"000000000000" when X = 283 AND Y = 61 else
"000000000000" when X = 284 AND Y = 61 else
"000000000000" when X = 285 AND Y = 61 else
"000000000000" when X = 286 AND Y = 61 else
"000000000000" when X = 287 AND Y = 61 else
"000000000000" when X = 288 AND Y = 61 else
"000000000000" when X = 289 AND Y = 61 else
"000000000000" when X = 290 AND Y = 61 else
"000000000000" when X = 291 AND Y = 61 else
"000000000000" when X = 292 AND Y = 61 else
"000000000000" when X = 293 AND Y = 61 else
"000000000000" when X = 294 AND Y = 61 else
"000000000000" when X = 295 AND Y = 61 else
"000000000000" when X = 296 AND Y = 61 else
"000000000000" when X = 297 AND Y = 61 else
"000000000000" when X = 298 AND Y = 61 else
"000000000000" when X = 299 AND Y = 61 else
"000000000000" when X = 300 AND Y = 61 else
"000000000000" when X = 301 AND Y = 61 else
"000000000000" when X = 302 AND Y = 61 else
"000000000000" when X = 303 AND Y = 61 else
"000000000000" when X = 304 AND Y = 61 else
"000000000000" when X = 305 AND Y = 61 else
"000000000000" when X = 306 AND Y = 61 else
"000000000000" when X = 307 AND Y = 61 else
"000000000000" when X = 308 AND Y = 61 else
"000000000000" when X = 309 AND Y = 61 else
"000000000000" when X = 310 AND Y = 61 else
"000000000000" when X = 311 AND Y = 61 else
"000000000000" when X = 312 AND Y = 61 else
"000000000000" when X = 313 AND Y = 61 else
"000000000000" when X = 314 AND Y = 61 else
"000000000000" when X = 315 AND Y = 61 else
"000000000000" when X = 316 AND Y = 61 else
"000000000000" when X = 317 AND Y = 61 else
"000000000000" when X = 318 AND Y = 61 else
"000000000000" when X = 319 AND Y = 61 else
"000000000000" when X = 320 AND Y = 61 else
"000000000000" when X = 321 AND Y = 61 else
"000000000000" when X = 322 AND Y = 61 else
"000000000000" when X = 323 AND Y = 61 else
"000000000000" when X = 324 AND Y = 61 else
"100010011101" when X = 0 AND Y = 62 else
"100010011101" when X = 1 AND Y = 62 else
"100010011101" when X = 2 AND Y = 62 else
"100010011101" when X = 3 AND Y = 62 else
"100010011101" when X = 4 AND Y = 62 else
"100010011101" when X = 5 AND Y = 62 else
"100010011101" when X = 6 AND Y = 62 else
"100010011101" when X = 7 AND Y = 62 else
"100010011101" when X = 8 AND Y = 62 else
"100010011101" when X = 9 AND Y = 62 else
"100010011101" when X = 10 AND Y = 62 else
"100010011101" when X = 11 AND Y = 62 else
"100010011101" when X = 12 AND Y = 62 else
"100010011101" when X = 13 AND Y = 62 else
"100010011101" when X = 14 AND Y = 62 else
"100010011101" when X = 15 AND Y = 62 else
"100010011101" when X = 16 AND Y = 62 else
"100010011101" when X = 17 AND Y = 62 else
"100010011101" when X = 18 AND Y = 62 else
"100010011101" when X = 19 AND Y = 62 else
"100010011101" when X = 20 AND Y = 62 else
"100010011101" when X = 21 AND Y = 62 else
"100010011101" when X = 22 AND Y = 62 else
"100010011101" when X = 23 AND Y = 62 else
"100010011101" when X = 24 AND Y = 62 else
"100010011101" when X = 25 AND Y = 62 else
"100010011101" when X = 26 AND Y = 62 else
"100010011101" when X = 27 AND Y = 62 else
"100010011101" when X = 28 AND Y = 62 else
"100010011101" when X = 29 AND Y = 62 else
"100010011101" when X = 30 AND Y = 62 else
"100010011101" when X = 31 AND Y = 62 else
"100010011101" when X = 32 AND Y = 62 else
"100010011101" when X = 33 AND Y = 62 else
"100010011101" when X = 34 AND Y = 62 else
"110111011111" when X = 35 AND Y = 62 else
"110111011111" when X = 36 AND Y = 62 else
"110111011111" when X = 37 AND Y = 62 else
"110111011111" when X = 38 AND Y = 62 else
"110111011111" when X = 39 AND Y = 62 else
"110111011111" when X = 40 AND Y = 62 else
"110111011111" when X = 41 AND Y = 62 else
"110111011111" when X = 42 AND Y = 62 else
"110111011111" when X = 43 AND Y = 62 else
"110111011111" when X = 44 AND Y = 62 else
"110111011111" when X = 45 AND Y = 62 else
"110111011111" when X = 46 AND Y = 62 else
"110111011111" when X = 47 AND Y = 62 else
"110111011111" when X = 48 AND Y = 62 else
"110111011111" when X = 49 AND Y = 62 else
"110111011111" when X = 50 AND Y = 62 else
"110111011111" when X = 51 AND Y = 62 else
"110111011111" when X = 52 AND Y = 62 else
"110111011111" when X = 53 AND Y = 62 else
"110111011111" when X = 54 AND Y = 62 else
"110111011111" when X = 55 AND Y = 62 else
"110111011111" when X = 56 AND Y = 62 else
"110111011111" when X = 57 AND Y = 62 else
"110111011111" when X = 58 AND Y = 62 else
"110111011111" when X = 59 AND Y = 62 else
"110111011111" when X = 60 AND Y = 62 else
"110111011111" when X = 61 AND Y = 62 else
"110111011111" when X = 62 AND Y = 62 else
"110111011111" when X = 63 AND Y = 62 else
"110111011111" when X = 64 AND Y = 62 else
"110111011111" when X = 65 AND Y = 62 else
"110111011111" when X = 66 AND Y = 62 else
"110111011111" when X = 67 AND Y = 62 else
"110111011111" when X = 68 AND Y = 62 else
"110111011111" when X = 69 AND Y = 62 else
"110111011111" when X = 70 AND Y = 62 else
"110111011111" when X = 71 AND Y = 62 else
"110111011111" when X = 72 AND Y = 62 else
"110111011111" when X = 73 AND Y = 62 else
"110111011111" when X = 74 AND Y = 62 else
"110111011111" when X = 75 AND Y = 62 else
"110111011111" when X = 76 AND Y = 62 else
"110111011111" when X = 77 AND Y = 62 else
"110111011111" when X = 78 AND Y = 62 else
"110111011111" when X = 79 AND Y = 62 else
"110111011111" when X = 80 AND Y = 62 else
"110111011111" when X = 81 AND Y = 62 else
"110111011111" when X = 82 AND Y = 62 else
"110111011111" when X = 83 AND Y = 62 else
"110111011111" when X = 84 AND Y = 62 else
"110111011111" when X = 85 AND Y = 62 else
"110111011111" when X = 86 AND Y = 62 else
"110111011111" when X = 87 AND Y = 62 else
"110111011111" when X = 88 AND Y = 62 else
"110111011111" when X = 89 AND Y = 62 else
"110111011111" when X = 90 AND Y = 62 else
"110111011111" when X = 91 AND Y = 62 else
"110111011111" when X = 92 AND Y = 62 else
"110111011111" when X = 93 AND Y = 62 else
"110111011111" when X = 94 AND Y = 62 else
"110111011111" when X = 95 AND Y = 62 else
"110111011111" when X = 96 AND Y = 62 else
"110111011111" when X = 97 AND Y = 62 else
"110111011111" when X = 98 AND Y = 62 else
"110111011111" when X = 99 AND Y = 62 else
"111111111111" when X = 100 AND Y = 62 else
"111111111111" when X = 101 AND Y = 62 else
"111111111111" when X = 102 AND Y = 62 else
"111111111111" when X = 103 AND Y = 62 else
"111111111111" when X = 104 AND Y = 62 else
"111111111111" when X = 105 AND Y = 62 else
"111111111111" when X = 106 AND Y = 62 else
"111111111111" when X = 107 AND Y = 62 else
"111111111111" when X = 108 AND Y = 62 else
"111111111111" when X = 109 AND Y = 62 else
"111111111111" when X = 110 AND Y = 62 else
"111111111111" when X = 111 AND Y = 62 else
"111111111111" when X = 112 AND Y = 62 else
"111111111111" when X = 113 AND Y = 62 else
"111111111111" when X = 114 AND Y = 62 else
"111111111111" when X = 115 AND Y = 62 else
"111111111111" when X = 116 AND Y = 62 else
"111111111111" when X = 117 AND Y = 62 else
"111111111111" when X = 118 AND Y = 62 else
"111111111111" when X = 119 AND Y = 62 else
"111111111111" when X = 120 AND Y = 62 else
"111111111111" when X = 121 AND Y = 62 else
"111111111111" when X = 122 AND Y = 62 else
"111111111111" when X = 123 AND Y = 62 else
"111111111111" when X = 124 AND Y = 62 else
"111111111111" when X = 125 AND Y = 62 else
"111111111111" when X = 126 AND Y = 62 else
"111111111111" when X = 127 AND Y = 62 else
"111111111111" when X = 128 AND Y = 62 else
"111111111111" when X = 129 AND Y = 62 else
"111111111111" when X = 130 AND Y = 62 else
"111111111111" when X = 131 AND Y = 62 else
"111111111111" when X = 132 AND Y = 62 else
"111111111111" when X = 133 AND Y = 62 else
"111111111111" when X = 134 AND Y = 62 else
"111111111111" when X = 135 AND Y = 62 else
"111111111111" when X = 136 AND Y = 62 else
"111111111111" when X = 137 AND Y = 62 else
"111111111111" when X = 138 AND Y = 62 else
"111111111111" when X = 139 AND Y = 62 else
"111111111111" when X = 140 AND Y = 62 else
"111111111111" when X = 141 AND Y = 62 else
"111111111111" when X = 142 AND Y = 62 else
"111111111111" when X = 143 AND Y = 62 else
"111111111111" when X = 144 AND Y = 62 else
"111111111111" when X = 145 AND Y = 62 else
"111111111111" when X = 146 AND Y = 62 else
"111111111111" when X = 147 AND Y = 62 else
"111111111111" when X = 148 AND Y = 62 else
"111111111111" when X = 149 AND Y = 62 else
"111111111111" when X = 150 AND Y = 62 else
"111111111111" when X = 151 AND Y = 62 else
"111111111111" when X = 152 AND Y = 62 else
"111111111111" when X = 153 AND Y = 62 else
"111111111111" when X = 154 AND Y = 62 else
"111111111111" when X = 155 AND Y = 62 else
"111111111111" when X = 156 AND Y = 62 else
"111111111111" when X = 157 AND Y = 62 else
"111111111111" when X = 158 AND Y = 62 else
"111111111111" when X = 159 AND Y = 62 else
"111111111111" when X = 160 AND Y = 62 else
"111111111111" when X = 161 AND Y = 62 else
"111111111111" when X = 162 AND Y = 62 else
"111111111111" when X = 163 AND Y = 62 else
"111111111111" when X = 164 AND Y = 62 else
"111111111111" when X = 165 AND Y = 62 else
"111111111111" when X = 166 AND Y = 62 else
"111111111111" when X = 167 AND Y = 62 else
"111111111111" when X = 168 AND Y = 62 else
"111111111111" when X = 169 AND Y = 62 else
"111111111111" when X = 170 AND Y = 62 else
"111111111111" when X = 171 AND Y = 62 else
"111111111111" when X = 172 AND Y = 62 else
"111111111111" when X = 173 AND Y = 62 else
"111111111111" when X = 174 AND Y = 62 else
"111111111111" when X = 175 AND Y = 62 else
"111111111111" when X = 176 AND Y = 62 else
"111111111111" when X = 177 AND Y = 62 else
"111111111111" when X = 178 AND Y = 62 else
"111111111111" when X = 179 AND Y = 62 else
"111111111111" when X = 180 AND Y = 62 else
"111111111111" when X = 181 AND Y = 62 else
"111111111111" when X = 182 AND Y = 62 else
"111111111111" when X = 183 AND Y = 62 else
"111111111111" when X = 184 AND Y = 62 else
"111111111111" when X = 185 AND Y = 62 else
"111111111111" when X = 186 AND Y = 62 else
"111111111111" when X = 187 AND Y = 62 else
"111111111111" when X = 188 AND Y = 62 else
"111111111111" when X = 189 AND Y = 62 else
"111111111111" when X = 190 AND Y = 62 else
"111111111111" when X = 191 AND Y = 62 else
"111111111111" when X = 192 AND Y = 62 else
"111111111111" when X = 193 AND Y = 62 else
"111111111111" when X = 194 AND Y = 62 else
"111111111111" when X = 195 AND Y = 62 else
"111111111111" when X = 196 AND Y = 62 else
"111111111111" when X = 197 AND Y = 62 else
"111111111111" when X = 198 AND Y = 62 else
"111111111111" when X = 199 AND Y = 62 else
"111111111111" when X = 200 AND Y = 62 else
"111111111111" when X = 201 AND Y = 62 else
"111111111111" when X = 202 AND Y = 62 else
"111111111111" when X = 203 AND Y = 62 else
"111111111111" when X = 204 AND Y = 62 else
"111111111111" when X = 205 AND Y = 62 else
"111111111111" when X = 206 AND Y = 62 else
"111111111111" when X = 207 AND Y = 62 else
"111111111111" when X = 208 AND Y = 62 else
"111111111111" when X = 209 AND Y = 62 else
"111111111111" when X = 210 AND Y = 62 else
"111111111111" when X = 211 AND Y = 62 else
"111111111111" when X = 212 AND Y = 62 else
"111111111111" when X = 213 AND Y = 62 else
"111111111111" when X = 214 AND Y = 62 else
"111111111111" when X = 215 AND Y = 62 else
"111111111111" when X = 216 AND Y = 62 else
"111111111111" when X = 217 AND Y = 62 else
"111111111111" when X = 218 AND Y = 62 else
"111111111111" when X = 219 AND Y = 62 else
"111111111111" when X = 220 AND Y = 62 else
"111111111111" when X = 221 AND Y = 62 else
"111111111111" when X = 222 AND Y = 62 else
"111111111111" when X = 223 AND Y = 62 else
"111111111111" when X = 224 AND Y = 62 else
"111111111111" when X = 225 AND Y = 62 else
"111111111111" when X = 226 AND Y = 62 else
"111111111111" when X = 227 AND Y = 62 else
"111111111111" when X = 228 AND Y = 62 else
"111111111111" when X = 229 AND Y = 62 else
"111111111111" when X = 230 AND Y = 62 else
"111111111111" when X = 231 AND Y = 62 else
"111111111111" when X = 232 AND Y = 62 else
"111111111111" when X = 233 AND Y = 62 else
"111111111111" when X = 234 AND Y = 62 else
"111111111111" when X = 235 AND Y = 62 else
"111111111111" when X = 236 AND Y = 62 else
"111111111111" when X = 237 AND Y = 62 else
"111111111111" when X = 238 AND Y = 62 else
"111111111111" when X = 239 AND Y = 62 else
"111111111111" when X = 240 AND Y = 62 else
"111111111111" when X = 241 AND Y = 62 else
"111111111111" when X = 242 AND Y = 62 else
"111111111111" when X = 243 AND Y = 62 else
"111111111111" when X = 244 AND Y = 62 else
"111111111111" when X = 245 AND Y = 62 else
"111111111111" when X = 246 AND Y = 62 else
"111111111111" when X = 247 AND Y = 62 else
"111111111111" when X = 248 AND Y = 62 else
"111111111111" when X = 249 AND Y = 62 else
"111111111111" when X = 250 AND Y = 62 else
"111111111111" when X = 251 AND Y = 62 else
"111111111111" when X = 252 AND Y = 62 else
"111111111111" when X = 253 AND Y = 62 else
"111111111111" when X = 254 AND Y = 62 else
"111111111111" when X = 255 AND Y = 62 else
"111111111111" when X = 256 AND Y = 62 else
"111111111111" when X = 257 AND Y = 62 else
"111111111111" when X = 258 AND Y = 62 else
"111111111111" when X = 259 AND Y = 62 else
"111111111111" when X = 260 AND Y = 62 else
"111111111111" when X = 261 AND Y = 62 else
"111111111111" when X = 262 AND Y = 62 else
"111111111111" when X = 263 AND Y = 62 else
"111111111111" when X = 264 AND Y = 62 else
"110111011111" when X = 265 AND Y = 62 else
"110111011111" when X = 266 AND Y = 62 else
"110111011111" when X = 267 AND Y = 62 else
"110111011111" when X = 268 AND Y = 62 else
"110111011111" when X = 269 AND Y = 62 else
"110111011111" when X = 270 AND Y = 62 else
"110111011111" when X = 271 AND Y = 62 else
"110111011111" when X = 272 AND Y = 62 else
"110111011111" when X = 273 AND Y = 62 else
"110111011111" when X = 274 AND Y = 62 else
"110111011111" when X = 275 AND Y = 62 else
"110111011111" when X = 276 AND Y = 62 else
"110111011111" when X = 277 AND Y = 62 else
"110111011111" when X = 278 AND Y = 62 else
"110111011111" when X = 279 AND Y = 62 else
"000000000000" when X = 280 AND Y = 62 else
"000000000000" when X = 281 AND Y = 62 else
"000000000000" when X = 282 AND Y = 62 else
"000000000000" when X = 283 AND Y = 62 else
"000000000000" when X = 284 AND Y = 62 else
"000000000000" when X = 285 AND Y = 62 else
"000000000000" when X = 286 AND Y = 62 else
"000000000000" when X = 287 AND Y = 62 else
"000000000000" when X = 288 AND Y = 62 else
"000000000000" when X = 289 AND Y = 62 else
"000000000000" when X = 290 AND Y = 62 else
"000000000000" when X = 291 AND Y = 62 else
"000000000000" when X = 292 AND Y = 62 else
"000000000000" when X = 293 AND Y = 62 else
"000000000000" when X = 294 AND Y = 62 else
"000000000000" when X = 295 AND Y = 62 else
"000000000000" when X = 296 AND Y = 62 else
"000000000000" when X = 297 AND Y = 62 else
"000000000000" when X = 298 AND Y = 62 else
"000000000000" when X = 299 AND Y = 62 else
"000000000000" when X = 300 AND Y = 62 else
"000000000000" when X = 301 AND Y = 62 else
"000000000000" when X = 302 AND Y = 62 else
"000000000000" when X = 303 AND Y = 62 else
"000000000000" when X = 304 AND Y = 62 else
"000000000000" when X = 305 AND Y = 62 else
"000000000000" when X = 306 AND Y = 62 else
"000000000000" when X = 307 AND Y = 62 else
"000000000000" when X = 308 AND Y = 62 else
"000000000000" when X = 309 AND Y = 62 else
"000000000000" when X = 310 AND Y = 62 else
"000000000000" when X = 311 AND Y = 62 else
"000000000000" when X = 312 AND Y = 62 else
"000000000000" when X = 313 AND Y = 62 else
"000000000000" when X = 314 AND Y = 62 else
"000000000000" when X = 315 AND Y = 62 else
"000000000000" when X = 316 AND Y = 62 else
"000000000000" when X = 317 AND Y = 62 else
"000000000000" when X = 318 AND Y = 62 else
"000000000000" when X = 319 AND Y = 62 else
"000000000000" when X = 320 AND Y = 62 else
"000000000000" when X = 321 AND Y = 62 else
"000000000000" when X = 322 AND Y = 62 else
"000000000000" when X = 323 AND Y = 62 else
"000000000000" when X = 324 AND Y = 62 else
"100010011101" when X = 0 AND Y = 63 else
"100010011101" when X = 1 AND Y = 63 else
"100010011101" when X = 2 AND Y = 63 else
"100010011101" when X = 3 AND Y = 63 else
"100010011101" when X = 4 AND Y = 63 else
"100010011101" when X = 5 AND Y = 63 else
"100010011101" when X = 6 AND Y = 63 else
"100010011101" when X = 7 AND Y = 63 else
"100010011101" when X = 8 AND Y = 63 else
"100010011101" when X = 9 AND Y = 63 else
"100010011101" when X = 10 AND Y = 63 else
"100010011101" when X = 11 AND Y = 63 else
"100010011101" when X = 12 AND Y = 63 else
"100010011101" when X = 13 AND Y = 63 else
"100010011101" when X = 14 AND Y = 63 else
"100010011101" when X = 15 AND Y = 63 else
"100010011101" when X = 16 AND Y = 63 else
"100010011101" when X = 17 AND Y = 63 else
"100010011101" when X = 18 AND Y = 63 else
"100010011101" when X = 19 AND Y = 63 else
"100010011101" when X = 20 AND Y = 63 else
"100010011101" when X = 21 AND Y = 63 else
"100010011101" when X = 22 AND Y = 63 else
"100010011101" when X = 23 AND Y = 63 else
"100010011101" when X = 24 AND Y = 63 else
"100010011101" when X = 25 AND Y = 63 else
"100010011101" when X = 26 AND Y = 63 else
"100010011101" when X = 27 AND Y = 63 else
"100010011101" when X = 28 AND Y = 63 else
"100010011101" when X = 29 AND Y = 63 else
"100010011101" when X = 30 AND Y = 63 else
"100010011101" when X = 31 AND Y = 63 else
"100010011101" when X = 32 AND Y = 63 else
"100010011101" when X = 33 AND Y = 63 else
"100010011101" when X = 34 AND Y = 63 else
"110111011111" when X = 35 AND Y = 63 else
"110111011111" when X = 36 AND Y = 63 else
"110111011111" when X = 37 AND Y = 63 else
"110111011111" when X = 38 AND Y = 63 else
"110111011111" when X = 39 AND Y = 63 else
"110111011111" when X = 40 AND Y = 63 else
"110111011111" when X = 41 AND Y = 63 else
"110111011111" when X = 42 AND Y = 63 else
"110111011111" when X = 43 AND Y = 63 else
"110111011111" when X = 44 AND Y = 63 else
"110111011111" when X = 45 AND Y = 63 else
"110111011111" when X = 46 AND Y = 63 else
"110111011111" when X = 47 AND Y = 63 else
"110111011111" when X = 48 AND Y = 63 else
"110111011111" when X = 49 AND Y = 63 else
"110111011111" when X = 50 AND Y = 63 else
"110111011111" when X = 51 AND Y = 63 else
"110111011111" when X = 52 AND Y = 63 else
"110111011111" when X = 53 AND Y = 63 else
"110111011111" when X = 54 AND Y = 63 else
"110111011111" when X = 55 AND Y = 63 else
"110111011111" when X = 56 AND Y = 63 else
"110111011111" when X = 57 AND Y = 63 else
"110111011111" when X = 58 AND Y = 63 else
"110111011111" when X = 59 AND Y = 63 else
"110111011111" when X = 60 AND Y = 63 else
"110111011111" when X = 61 AND Y = 63 else
"110111011111" when X = 62 AND Y = 63 else
"110111011111" when X = 63 AND Y = 63 else
"110111011111" when X = 64 AND Y = 63 else
"110111011111" when X = 65 AND Y = 63 else
"110111011111" when X = 66 AND Y = 63 else
"110111011111" when X = 67 AND Y = 63 else
"110111011111" when X = 68 AND Y = 63 else
"110111011111" when X = 69 AND Y = 63 else
"110111011111" when X = 70 AND Y = 63 else
"110111011111" when X = 71 AND Y = 63 else
"110111011111" when X = 72 AND Y = 63 else
"110111011111" when X = 73 AND Y = 63 else
"110111011111" when X = 74 AND Y = 63 else
"110111011111" when X = 75 AND Y = 63 else
"110111011111" when X = 76 AND Y = 63 else
"110111011111" when X = 77 AND Y = 63 else
"110111011111" when X = 78 AND Y = 63 else
"110111011111" when X = 79 AND Y = 63 else
"110111011111" when X = 80 AND Y = 63 else
"110111011111" when X = 81 AND Y = 63 else
"110111011111" when X = 82 AND Y = 63 else
"110111011111" when X = 83 AND Y = 63 else
"110111011111" when X = 84 AND Y = 63 else
"110111011111" when X = 85 AND Y = 63 else
"110111011111" when X = 86 AND Y = 63 else
"110111011111" when X = 87 AND Y = 63 else
"110111011111" when X = 88 AND Y = 63 else
"110111011111" when X = 89 AND Y = 63 else
"110111011111" when X = 90 AND Y = 63 else
"110111011111" when X = 91 AND Y = 63 else
"110111011111" when X = 92 AND Y = 63 else
"110111011111" when X = 93 AND Y = 63 else
"110111011111" when X = 94 AND Y = 63 else
"110111011111" when X = 95 AND Y = 63 else
"110111011111" when X = 96 AND Y = 63 else
"110111011111" when X = 97 AND Y = 63 else
"110111011111" when X = 98 AND Y = 63 else
"110111011111" when X = 99 AND Y = 63 else
"111111111111" when X = 100 AND Y = 63 else
"111111111111" when X = 101 AND Y = 63 else
"111111111111" when X = 102 AND Y = 63 else
"111111111111" when X = 103 AND Y = 63 else
"111111111111" when X = 104 AND Y = 63 else
"111111111111" when X = 105 AND Y = 63 else
"111111111111" when X = 106 AND Y = 63 else
"111111111111" when X = 107 AND Y = 63 else
"111111111111" when X = 108 AND Y = 63 else
"111111111111" when X = 109 AND Y = 63 else
"111111111111" when X = 110 AND Y = 63 else
"111111111111" when X = 111 AND Y = 63 else
"111111111111" when X = 112 AND Y = 63 else
"111111111111" when X = 113 AND Y = 63 else
"111111111111" when X = 114 AND Y = 63 else
"111111111111" when X = 115 AND Y = 63 else
"111111111111" when X = 116 AND Y = 63 else
"111111111111" when X = 117 AND Y = 63 else
"111111111111" when X = 118 AND Y = 63 else
"111111111111" when X = 119 AND Y = 63 else
"111111111111" when X = 120 AND Y = 63 else
"111111111111" when X = 121 AND Y = 63 else
"111111111111" when X = 122 AND Y = 63 else
"111111111111" when X = 123 AND Y = 63 else
"111111111111" when X = 124 AND Y = 63 else
"111111111111" when X = 125 AND Y = 63 else
"111111111111" when X = 126 AND Y = 63 else
"111111111111" when X = 127 AND Y = 63 else
"111111111111" when X = 128 AND Y = 63 else
"111111111111" when X = 129 AND Y = 63 else
"111111111111" when X = 130 AND Y = 63 else
"111111111111" when X = 131 AND Y = 63 else
"111111111111" when X = 132 AND Y = 63 else
"111111111111" when X = 133 AND Y = 63 else
"111111111111" when X = 134 AND Y = 63 else
"111111111111" when X = 135 AND Y = 63 else
"111111111111" when X = 136 AND Y = 63 else
"111111111111" when X = 137 AND Y = 63 else
"111111111111" when X = 138 AND Y = 63 else
"111111111111" when X = 139 AND Y = 63 else
"111111111111" when X = 140 AND Y = 63 else
"111111111111" when X = 141 AND Y = 63 else
"111111111111" when X = 142 AND Y = 63 else
"111111111111" when X = 143 AND Y = 63 else
"111111111111" when X = 144 AND Y = 63 else
"111111111111" when X = 145 AND Y = 63 else
"111111111111" when X = 146 AND Y = 63 else
"111111111111" when X = 147 AND Y = 63 else
"111111111111" when X = 148 AND Y = 63 else
"111111111111" when X = 149 AND Y = 63 else
"111111111111" when X = 150 AND Y = 63 else
"111111111111" when X = 151 AND Y = 63 else
"111111111111" when X = 152 AND Y = 63 else
"111111111111" when X = 153 AND Y = 63 else
"111111111111" when X = 154 AND Y = 63 else
"111111111111" when X = 155 AND Y = 63 else
"111111111111" when X = 156 AND Y = 63 else
"111111111111" when X = 157 AND Y = 63 else
"111111111111" when X = 158 AND Y = 63 else
"111111111111" when X = 159 AND Y = 63 else
"111111111111" when X = 160 AND Y = 63 else
"111111111111" when X = 161 AND Y = 63 else
"111111111111" when X = 162 AND Y = 63 else
"111111111111" when X = 163 AND Y = 63 else
"111111111111" when X = 164 AND Y = 63 else
"111111111111" when X = 165 AND Y = 63 else
"111111111111" when X = 166 AND Y = 63 else
"111111111111" when X = 167 AND Y = 63 else
"111111111111" when X = 168 AND Y = 63 else
"111111111111" when X = 169 AND Y = 63 else
"111111111111" when X = 170 AND Y = 63 else
"111111111111" when X = 171 AND Y = 63 else
"111111111111" when X = 172 AND Y = 63 else
"111111111111" when X = 173 AND Y = 63 else
"111111111111" when X = 174 AND Y = 63 else
"111111111111" when X = 175 AND Y = 63 else
"111111111111" when X = 176 AND Y = 63 else
"111111111111" when X = 177 AND Y = 63 else
"111111111111" when X = 178 AND Y = 63 else
"111111111111" when X = 179 AND Y = 63 else
"111111111111" when X = 180 AND Y = 63 else
"111111111111" when X = 181 AND Y = 63 else
"111111111111" when X = 182 AND Y = 63 else
"111111111111" when X = 183 AND Y = 63 else
"111111111111" when X = 184 AND Y = 63 else
"111111111111" when X = 185 AND Y = 63 else
"111111111111" when X = 186 AND Y = 63 else
"111111111111" when X = 187 AND Y = 63 else
"111111111111" when X = 188 AND Y = 63 else
"111111111111" when X = 189 AND Y = 63 else
"111111111111" when X = 190 AND Y = 63 else
"111111111111" when X = 191 AND Y = 63 else
"111111111111" when X = 192 AND Y = 63 else
"111111111111" when X = 193 AND Y = 63 else
"111111111111" when X = 194 AND Y = 63 else
"111111111111" when X = 195 AND Y = 63 else
"111111111111" when X = 196 AND Y = 63 else
"111111111111" when X = 197 AND Y = 63 else
"111111111111" when X = 198 AND Y = 63 else
"111111111111" when X = 199 AND Y = 63 else
"111111111111" when X = 200 AND Y = 63 else
"111111111111" when X = 201 AND Y = 63 else
"111111111111" when X = 202 AND Y = 63 else
"111111111111" when X = 203 AND Y = 63 else
"111111111111" when X = 204 AND Y = 63 else
"111111111111" when X = 205 AND Y = 63 else
"111111111111" when X = 206 AND Y = 63 else
"111111111111" when X = 207 AND Y = 63 else
"111111111111" when X = 208 AND Y = 63 else
"111111111111" when X = 209 AND Y = 63 else
"111111111111" when X = 210 AND Y = 63 else
"111111111111" when X = 211 AND Y = 63 else
"111111111111" when X = 212 AND Y = 63 else
"111111111111" when X = 213 AND Y = 63 else
"111111111111" when X = 214 AND Y = 63 else
"111111111111" when X = 215 AND Y = 63 else
"111111111111" when X = 216 AND Y = 63 else
"111111111111" when X = 217 AND Y = 63 else
"111111111111" when X = 218 AND Y = 63 else
"111111111111" when X = 219 AND Y = 63 else
"111111111111" when X = 220 AND Y = 63 else
"111111111111" when X = 221 AND Y = 63 else
"111111111111" when X = 222 AND Y = 63 else
"111111111111" when X = 223 AND Y = 63 else
"111111111111" when X = 224 AND Y = 63 else
"111111111111" when X = 225 AND Y = 63 else
"111111111111" when X = 226 AND Y = 63 else
"111111111111" when X = 227 AND Y = 63 else
"111111111111" when X = 228 AND Y = 63 else
"111111111111" when X = 229 AND Y = 63 else
"111111111111" when X = 230 AND Y = 63 else
"111111111111" when X = 231 AND Y = 63 else
"111111111111" when X = 232 AND Y = 63 else
"111111111111" when X = 233 AND Y = 63 else
"111111111111" when X = 234 AND Y = 63 else
"111111111111" when X = 235 AND Y = 63 else
"111111111111" when X = 236 AND Y = 63 else
"111111111111" when X = 237 AND Y = 63 else
"111111111111" when X = 238 AND Y = 63 else
"111111111111" when X = 239 AND Y = 63 else
"111111111111" when X = 240 AND Y = 63 else
"111111111111" when X = 241 AND Y = 63 else
"111111111111" when X = 242 AND Y = 63 else
"111111111111" when X = 243 AND Y = 63 else
"111111111111" when X = 244 AND Y = 63 else
"111111111111" when X = 245 AND Y = 63 else
"111111111111" when X = 246 AND Y = 63 else
"111111111111" when X = 247 AND Y = 63 else
"111111111111" when X = 248 AND Y = 63 else
"111111111111" when X = 249 AND Y = 63 else
"111111111111" when X = 250 AND Y = 63 else
"111111111111" when X = 251 AND Y = 63 else
"111111111111" when X = 252 AND Y = 63 else
"111111111111" when X = 253 AND Y = 63 else
"111111111111" when X = 254 AND Y = 63 else
"111111111111" when X = 255 AND Y = 63 else
"111111111111" when X = 256 AND Y = 63 else
"111111111111" when X = 257 AND Y = 63 else
"111111111111" when X = 258 AND Y = 63 else
"111111111111" when X = 259 AND Y = 63 else
"111111111111" when X = 260 AND Y = 63 else
"111111111111" when X = 261 AND Y = 63 else
"111111111111" when X = 262 AND Y = 63 else
"111111111111" when X = 263 AND Y = 63 else
"111111111111" when X = 264 AND Y = 63 else
"110111011111" when X = 265 AND Y = 63 else
"110111011111" when X = 266 AND Y = 63 else
"110111011111" when X = 267 AND Y = 63 else
"110111011111" when X = 268 AND Y = 63 else
"110111011111" when X = 269 AND Y = 63 else
"110111011111" when X = 270 AND Y = 63 else
"110111011111" when X = 271 AND Y = 63 else
"110111011111" when X = 272 AND Y = 63 else
"110111011111" when X = 273 AND Y = 63 else
"110111011111" when X = 274 AND Y = 63 else
"110111011111" when X = 275 AND Y = 63 else
"110111011111" when X = 276 AND Y = 63 else
"110111011111" when X = 277 AND Y = 63 else
"110111011111" when X = 278 AND Y = 63 else
"110111011111" when X = 279 AND Y = 63 else
"000000000000" when X = 280 AND Y = 63 else
"000000000000" when X = 281 AND Y = 63 else
"000000000000" when X = 282 AND Y = 63 else
"000000000000" when X = 283 AND Y = 63 else
"000000000000" when X = 284 AND Y = 63 else
"000000000000" when X = 285 AND Y = 63 else
"000000000000" when X = 286 AND Y = 63 else
"000000000000" when X = 287 AND Y = 63 else
"000000000000" when X = 288 AND Y = 63 else
"000000000000" when X = 289 AND Y = 63 else
"000000000000" when X = 290 AND Y = 63 else
"000000000000" when X = 291 AND Y = 63 else
"000000000000" when X = 292 AND Y = 63 else
"000000000000" when X = 293 AND Y = 63 else
"000000000000" when X = 294 AND Y = 63 else
"000000000000" when X = 295 AND Y = 63 else
"000000000000" when X = 296 AND Y = 63 else
"000000000000" when X = 297 AND Y = 63 else
"000000000000" when X = 298 AND Y = 63 else
"000000000000" when X = 299 AND Y = 63 else
"000000000000" when X = 300 AND Y = 63 else
"000000000000" when X = 301 AND Y = 63 else
"000000000000" when X = 302 AND Y = 63 else
"000000000000" when X = 303 AND Y = 63 else
"000000000000" when X = 304 AND Y = 63 else
"000000000000" when X = 305 AND Y = 63 else
"000000000000" when X = 306 AND Y = 63 else
"000000000000" when X = 307 AND Y = 63 else
"000000000000" when X = 308 AND Y = 63 else
"000000000000" when X = 309 AND Y = 63 else
"000000000000" when X = 310 AND Y = 63 else
"000000000000" when X = 311 AND Y = 63 else
"000000000000" when X = 312 AND Y = 63 else
"000000000000" when X = 313 AND Y = 63 else
"000000000000" when X = 314 AND Y = 63 else
"000000000000" when X = 315 AND Y = 63 else
"000000000000" when X = 316 AND Y = 63 else
"000000000000" when X = 317 AND Y = 63 else
"000000000000" when X = 318 AND Y = 63 else
"000000000000" when X = 319 AND Y = 63 else
"000000000000" when X = 320 AND Y = 63 else
"000000000000" when X = 321 AND Y = 63 else
"000000000000" when X = 322 AND Y = 63 else
"000000000000" when X = 323 AND Y = 63 else
"000000000000" when X = 324 AND Y = 63 else
"100010011101" when X = 0 AND Y = 64 else
"100010011101" when X = 1 AND Y = 64 else
"100010011101" when X = 2 AND Y = 64 else
"100010011101" when X = 3 AND Y = 64 else
"100010011101" when X = 4 AND Y = 64 else
"100010011101" when X = 5 AND Y = 64 else
"100010011101" when X = 6 AND Y = 64 else
"100010011101" when X = 7 AND Y = 64 else
"100010011101" when X = 8 AND Y = 64 else
"100010011101" when X = 9 AND Y = 64 else
"100010011101" when X = 10 AND Y = 64 else
"100010011101" when X = 11 AND Y = 64 else
"100010011101" when X = 12 AND Y = 64 else
"100010011101" when X = 13 AND Y = 64 else
"100010011101" when X = 14 AND Y = 64 else
"100010011101" when X = 15 AND Y = 64 else
"100010011101" when X = 16 AND Y = 64 else
"100010011101" when X = 17 AND Y = 64 else
"100010011101" when X = 18 AND Y = 64 else
"100010011101" when X = 19 AND Y = 64 else
"100010011101" when X = 20 AND Y = 64 else
"100010011101" when X = 21 AND Y = 64 else
"100010011101" when X = 22 AND Y = 64 else
"100010011101" when X = 23 AND Y = 64 else
"100010011101" when X = 24 AND Y = 64 else
"100010011101" when X = 25 AND Y = 64 else
"100010011101" when X = 26 AND Y = 64 else
"100010011101" when X = 27 AND Y = 64 else
"100010011101" when X = 28 AND Y = 64 else
"100010011101" when X = 29 AND Y = 64 else
"100010011101" when X = 30 AND Y = 64 else
"100010011101" when X = 31 AND Y = 64 else
"100010011101" when X = 32 AND Y = 64 else
"100010011101" when X = 33 AND Y = 64 else
"100010011101" when X = 34 AND Y = 64 else
"110111011111" when X = 35 AND Y = 64 else
"110111011111" when X = 36 AND Y = 64 else
"110111011111" when X = 37 AND Y = 64 else
"110111011111" when X = 38 AND Y = 64 else
"110111011111" when X = 39 AND Y = 64 else
"110111011111" when X = 40 AND Y = 64 else
"110111011111" when X = 41 AND Y = 64 else
"110111011111" when X = 42 AND Y = 64 else
"110111011111" when X = 43 AND Y = 64 else
"110111011111" when X = 44 AND Y = 64 else
"110111011111" when X = 45 AND Y = 64 else
"110111011111" when X = 46 AND Y = 64 else
"110111011111" when X = 47 AND Y = 64 else
"110111011111" when X = 48 AND Y = 64 else
"110111011111" when X = 49 AND Y = 64 else
"110111011111" when X = 50 AND Y = 64 else
"110111011111" when X = 51 AND Y = 64 else
"110111011111" when X = 52 AND Y = 64 else
"110111011111" when X = 53 AND Y = 64 else
"110111011111" when X = 54 AND Y = 64 else
"110111011111" when X = 55 AND Y = 64 else
"110111011111" when X = 56 AND Y = 64 else
"110111011111" when X = 57 AND Y = 64 else
"110111011111" when X = 58 AND Y = 64 else
"110111011111" when X = 59 AND Y = 64 else
"110111011111" when X = 60 AND Y = 64 else
"110111011111" when X = 61 AND Y = 64 else
"110111011111" when X = 62 AND Y = 64 else
"110111011111" when X = 63 AND Y = 64 else
"110111011111" when X = 64 AND Y = 64 else
"110111011111" when X = 65 AND Y = 64 else
"110111011111" when X = 66 AND Y = 64 else
"110111011111" when X = 67 AND Y = 64 else
"110111011111" when X = 68 AND Y = 64 else
"110111011111" when X = 69 AND Y = 64 else
"110111011111" when X = 70 AND Y = 64 else
"110111011111" when X = 71 AND Y = 64 else
"110111011111" when X = 72 AND Y = 64 else
"110111011111" when X = 73 AND Y = 64 else
"110111011111" when X = 74 AND Y = 64 else
"110111011111" when X = 75 AND Y = 64 else
"110111011111" when X = 76 AND Y = 64 else
"110111011111" when X = 77 AND Y = 64 else
"110111011111" when X = 78 AND Y = 64 else
"110111011111" when X = 79 AND Y = 64 else
"110111011111" when X = 80 AND Y = 64 else
"110111011111" when X = 81 AND Y = 64 else
"110111011111" when X = 82 AND Y = 64 else
"110111011111" when X = 83 AND Y = 64 else
"110111011111" when X = 84 AND Y = 64 else
"110111011111" when X = 85 AND Y = 64 else
"110111011111" when X = 86 AND Y = 64 else
"110111011111" when X = 87 AND Y = 64 else
"110111011111" when X = 88 AND Y = 64 else
"110111011111" when X = 89 AND Y = 64 else
"110111011111" when X = 90 AND Y = 64 else
"110111011111" when X = 91 AND Y = 64 else
"110111011111" when X = 92 AND Y = 64 else
"110111011111" when X = 93 AND Y = 64 else
"110111011111" when X = 94 AND Y = 64 else
"110111011111" when X = 95 AND Y = 64 else
"110111011111" when X = 96 AND Y = 64 else
"110111011111" when X = 97 AND Y = 64 else
"110111011111" when X = 98 AND Y = 64 else
"110111011111" when X = 99 AND Y = 64 else
"111111111111" when X = 100 AND Y = 64 else
"111111111111" when X = 101 AND Y = 64 else
"111111111111" when X = 102 AND Y = 64 else
"111111111111" when X = 103 AND Y = 64 else
"111111111111" when X = 104 AND Y = 64 else
"111111111111" when X = 105 AND Y = 64 else
"111111111111" when X = 106 AND Y = 64 else
"111111111111" when X = 107 AND Y = 64 else
"111111111111" when X = 108 AND Y = 64 else
"111111111111" when X = 109 AND Y = 64 else
"111111111111" when X = 110 AND Y = 64 else
"111111111111" when X = 111 AND Y = 64 else
"111111111111" when X = 112 AND Y = 64 else
"111111111111" when X = 113 AND Y = 64 else
"111111111111" when X = 114 AND Y = 64 else
"111111111111" when X = 115 AND Y = 64 else
"111111111111" when X = 116 AND Y = 64 else
"111111111111" when X = 117 AND Y = 64 else
"111111111111" when X = 118 AND Y = 64 else
"111111111111" when X = 119 AND Y = 64 else
"111111111111" when X = 120 AND Y = 64 else
"111111111111" when X = 121 AND Y = 64 else
"111111111111" when X = 122 AND Y = 64 else
"111111111111" when X = 123 AND Y = 64 else
"111111111111" when X = 124 AND Y = 64 else
"111111111111" when X = 125 AND Y = 64 else
"111111111111" when X = 126 AND Y = 64 else
"111111111111" when X = 127 AND Y = 64 else
"111111111111" when X = 128 AND Y = 64 else
"111111111111" when X = 129 AND Y = 64 else
"111111111111" when X = 130 AND Y = 64 else
"111111111111" when X = 131 AND Y = 64 else
"111111111111" when X = 132 AND Y = 64 else
"111111111111" when X = 133 AND Y = 64 else
"111111111111" when X = 134 AND Y = 64 else
"111111111111" when X = 135 AND Y = 64 else
"111111111111" when X = 136 AND Y = 64 else
"111111111111" when X = 137 AND Y = 64 else
"111111111111" when X = 138 AND Y = 64 else
"111111111111" when X = 139 AND Y = 64 else
"111111111111" when X = 140 AND Y = 64 else
"111111111111" when X = 141 AND Y = 64 else
"111111111111" when X = 142 AND Y = 64 else
"111111111111" when X = 143 AND Y = 64 else
"111111111111" when X = 144 AND Y = 64 else
"111111111111" when X = 145 AND Y = 64 else
"111111111111" when X = 146 AND Y = 64 else
"111111111111" when X = 147 AND Y = 64 else
"111111111111" when X = 148 AND Y = 64 else
"111111111111" when X = 149 AND Y = 64 else
"111111111111" when X = 150 AND Y = 64 else
"111111111111" when X = 151 AND Y = 64 else
"111111111111" when X = 152 AND Y = 64 else
"111111111111" when X = 153 AND Y = 64 else
"111111111111" when X = 154 AND Y = 64 else
"111111111111" when X = 155 AND Y = 64 else
"111111111111" when X = 156 AND Y = 64 else
"111111111111" when X = 157 AND Y = 64 else
"111111111111" when X = 158 AND Y = 64 else
"111111111111" when X = 159 AND Y = 64 else
"111111111111" when X = 160 AND Y = 64 else
"111111111111" when X = 161 AND Y = 64 else
"111111111111" when X = 162 AND Y = 64 else
"111111111111" when X = 163 AND Y = 64 else
"111111111111" when X = 164 AND Y = 64 else
"111111111111" when X = 165 AND Y = 64 else
"111111111111" when X = 166 AND Y = 64 else
"111111111111" when X = 167 AND Y = 64 else
"111111111111" when X = 168 AND Y = 64 else
"111111111111" when X = 169 AND Y = 64 else
"111111111111" when X = 170 AND Y = 64 else
"111111111111" when X = 171 AND Y = 64 else
"111111111111" when X = 172 AND Y = 64 else
"111111111111" when X = 173 AND Y = 64 else
"111111111111" when X = 174 AND Y = 64 else
"111111111111" when X = 175 AND Y = 64 else
"111111111111" when X = 176 AND Y = 64 else
"111111111111" when X = 177 AND Y = 64 else
"111111111111" when X = 178 AND Y = 64 else
"111111111111" when X = 179 AND Y = 64 else
"111111111111" when X = 180 AND Y = 64 else
"111111111111" when X = 181 AND Y = 64 else
"111111111111" when X = 182 AND Y = 64 else
"111111111111" when X = 183 AND Y = 64 else
"111111111111" when X = 184 AND Y = 64 else
"111111111111" when X = 185 AND Y = 64 else
"111111111111" when X = 186 AND Y = 64 else
"111111111111" when X = 187 AND Y = 64 else
"111111111111" when X = 188 AND Y = 64 else
"111111111111" when X = 189 AND Y = 64 else
"111111111111" when X = 190 AND Y = 64 else
"111111111111" when X = 191 AND Y = 64 else
"111111111111" when X = 192 AND Y = 64 else
"111111111111" when X = 193 AND Y = 64 else
"111111111111" when X = 194 AND Y = 64 else
"111111111111" when X = 195 AND Y = 64 else
"111111111111" when X = 196 AND Y = 64 else
"111111111111" when X = 197 AND Y = 64 else
"111111111111" when X = 198 AND Y = 64 else
"111111111111" when X = 199 AND Y = 64 else
"111111111111" when X = 200 AND Y = 64 else
"111111111111" when X = 201 AND Y = 64 else
"111111111111" when X = 202 AND Y = 64 else
"111111111111" when X = 203 AND Y = 64 else
"111111111111" when X = 204 AND Y = 64 else
"111111111111" when X = 205 AND Y = 64 else
"111111111111" when X = 206 AND Y = 64 else
"111111111111" when X = 207 AND Y = 64 else
"111111111111" when X = 208 AND Y = 64 else
"111111111111" when X = 209 AND Y = 64 else
"111111111111" when X = 210 AND Y = 64 else
"111111111111" when X = 211 AND Y = 64 else
"111111111111" when X = 212 AND Y = 64 else
"111111111111" when X = 213 AND Y = 64 else
"111111111111" when X = 214 AND Y = 64 else
"111111111111" when X = 215 AND Y = 64 else
"111111111111" when X = 216 AND Y = 64 else
"111111111111" when X = 217 AND Y = 64 else
"111111111111" when X = 218 AND Y = 64 else
"111111111111" when X = 219 AND Y = 64 else
"111111111111" when X = 220 AND Y = 64 else
"111111111111" when X = 221 AND Y = 64 else
"111111111111" when X = 222 AND Y = 64 else
"111111111111" when X = 223 AND Y = 64 else
"111111111111" when X = 224 AND Y = 64 else
"111111111111" when X = 225 AND Y = 64 else
"111111111111" when X = 226 AND Y = 64 else
"111111111111" when X = 227 AND Y = 64 else
"111111111111" when X = 228 AND Y = 64 else
"111111111111" when X = 229 AND Y = 64 else
"111111111111" when X = 230 AND Y = 64 else
"111111111111" when X = 231 AND Y = 64 else
"111111111111" when X = 232 AND Y = 64 else
"111111111111" when X = 233 AND Y = 64 else
"111111111111" when X = 234 AND Y = 64 else
"111111111111" when X = 235 AND Y = 64 else
"111111111111" when X = 236 AND Y = 64 else
"111111111111" when X = 237 AND Y = 64 else
"111111111111" when X = 238 AND Y = 64 else
"111111111111" when X = 239 AND Y = 64 else
"111111111111" when X = 240 AND Y = 64 else
"111111111111" when X = 241 AND Y = 64 else
"111111111111" when X = 242 AND Y = 64 else
"111111111111" when X = 243 AND Y = 64 else
"111111111111" when X = 244 AND Y = 64 else
"111111111111" when X = 245 AND Y = 64 else
"111111111111" when X = 246 AND Y = 64 else
"111111111111" when X = 247 AND Y = 64 else
"111111111111" when X = 248 AND Y = 64 else
"111111111111" when X = 249 AND Y = 64 else
"111111111111" when X = 250 AND Y = 64 else
"111111111111" when X = 251 AND Y = 64 else
"111111111111" when X = 252 AND Y = 64 else
"111111111111" when X = 253 AND Y = 64 else
"111111111111" when X = 254 AND Y = 64 else
"111111111111" when X = 255 AND Y = 64 else
"111111111111" when X = 256 AND Y = 64 else
"111111111111" when X = 257 AND Y = 64 else
"111111111111" when X = 258 AND Y = 64 else
"111111111111" when X = 259 AND Y = 64 else
"111111111111" when X = 260 AND Y = 64 else
"111111111111" when X = 261 AND Y = 64 else
"111111111111" when X = 262 AND Y = 64 else
"111111111111" when X = 263 AND Y = 64 else
"111111111111" when X = 264 AND Y = 64 else
"110111011111" when X = 265 AND Y = 64 else
"110111011111" when X = 266 AND Y = 64 else
"110111011111" when X = 267 AND Y = 64 else
"110111011111" when X = 268 AND Y = 64 else
"110111011111" when X = 269 AND Y = 64 else
"110111011111" when X = 270 AND Y = 64 else
"110111011111" when X = 271 AND Y = 64 else
"110111011111" when X = 272 AND Y = 64 else
"110111011111" when X = 273 AND Y = 64 else
"110111011111" when X = 274 AND Y = 64 else
"110111011111" when X = 275 AND Y = 64 else
"110111011111" when X = 276 AND Y = 64 else
"110111011111" when X = 277 AND Y = 64 else
"110111011111" when X = 278 AND Y = 64 else
"110111011111" when X = 279 AND Y = 64 else
"000000000000" when X = 280 AND Y = 64 else
"000000000000" when X = 281 AND Y = 64 else
"000000000000" when X = 282 AND Y = 64 else
"000000000000" when X = 283 AND Y = 64 else
"000000000000" when X = 284 AND Y = 64 else
"000000000000" when X = 285 AND Y = 64 else
"000000000000" when X = 286 AND Y = 64 else
"000000000000" when X = 287 AND Y = 64 else
"000000000000" when X = 288 AND Y = 64 else
"000000000000" when X = 289 AND Y = 64 else
"000000000000" when X = 290 AND Y = 64 else
"000000000000" when X = 291 AND Y = 64 else
"000000000000" when X = 292 AND Y = 64 else
"000000000000" when X = 293 AND Y = 64 else
"000000000000" when X = 294 AND Y = 64 else
"000000000000" when X = 295 AND Y = 64 else
"000000000000" when X = 296 AND Y = 64 else
"000000000000" when X = 297 AND Y = 64 else
"000000000000" when X = 298 AND Y = 64 else
"000000000000" when X = 299 AND Y = 64 else
"000000000000" when X = 300 AND Y = 64 else
"000000000000" when X = 301 AND Y = 64 else
"000000000000" when X = 302 AND Y = 64 else
"000000000000" when X = 303 AND Y = 64 else
"000000000000" when X = 304 AND Y = 64 else
"000000000000" when X = 305 AND Y = 64 else
"000000000000" when X = 306 AND Y = 64 else
"000000000000" when X = 307 AND Y = 64 else
"000000000000" when X = 308 AND Y = 64 else
"000000000000" when X = 309 AND Y = 64 else
"000000000000" when X = 310 AND Y = 64 else
"000000000000" when X = 311 AND Y = 64 else
"000000000000" when X = 312 AND Y = 64 else
"000000000000" when X = 313 AND Y = 64 else
"000000000000" when X = 314 AND Y = 64 else
"000000000000" when X = 315 AND Y = 64 else
"000000000000" when X = 316 AND Y = 64 else
"000000000000" when X = 317 AND Y = 64 else
"000000000000" when X = 318 AND Y = 64 else
"000000000000" when X = 319 AND Y = 64 else
"000000000000" when X = 320 AND Y = 64 else
"000000000000" when X = 321 AND Y = 64 else
"000000000000" when X = 322 AND Y = 64 else
"000000000000" when X = 323 AND Y = 64 else
"000000000000" when X = 324 AND Y = 64 else
"100010011101" when X = 0 AND Y = 65 else
"100010011101" when X = 1 AND Y = 65 else
"100010011101" when X = 2 AND Y = 65 else
"100010011101" when X = 3 AND Y = 65 else
"100010011101" when X = 4 AND Y = 65 else
"100010011101" when X = 5 AND Y = 65 else
"100010011101" when X = 6 AND Y = 65 else
"100010011101" when X = 7 AND Y = 65 else
"100010011101" when X = 8 AND Y = 65 else
"100010011101" when X = 9 AND Y = 65 else
"100010011101" when X = 10 AND Y = 65 else
"100010011101" when X = 11 AND Y = 65 else
"100010011101" when X = 12 AND Y = 65 else
"100010011101" when X = 13 AND Y = 65 else
"100010011101" when X = 14 AND Y = 65 else
"100010011101" when X = 15 AND Y = 65 else
"100010011101" when X = 16 AND Y = 65 else
"100010011101" when X = 17 AND Y = 65 else
"100010011101" when X = 18 AND Y = 65 else
"100010011101" when X = 19 AND Y = 65 else
"100010011101" when X = 20 AND Y = 65 else
"100010011101" when X = 21 AND Y = 65 else
"100010011101" when X = 22 AND Y = 65 else
"100010011101" when X = 23 AND Y = 65 else
"100010011101" when X = 24 AND Y = 65 else
"100010011101" when X = 25 AND Y = 65 else
"100010011101" when X = 26 AND Y = 65 else
"100010011101" when X = 27 AND Y = 65 else
"100010011101" when X = 28 AND Y = 65 else
"100010011101" when X = 29 AND Y = 65 else
"100010011101" when X = 30 AND Y = 65 else
"100010011101" when X = 31 AND Y = 65 else
"100010011101" when X = 32 AND Y = 65 else
"100010011101" when X = 33 AND Y = 65 else
"100010011101" when X = 34 AND Y = 65 else
"110111011111" when X = 35 AND Y = 65 else
"110111011111" when X = 36 AND Y = 65 else
"110111011111" when X = 37 AND Y = 65 else
"110111011111" when X = 38 AND Y = 65 else
"110111011111" when X = 39 AND Y = 65 else
"110111011111" when X = 40 AND Y = 65 else
"110111011111" when X = 41 AND Y = 65 else
"110111011111" when X = 42 AND Y = 65 else
"110111011111" when X = 43 AND Y = 65 else
"110111011111" when X = 44 AND Y = 65 else
"110111011111" when X = 45 AND Y = 65 else
"110111011111" when X = 46 AND Y = 65 else
"110111011111" when X = 47 AND Y = 65 else
"110111011111" when X = 48 AND Y = 65 else
"110111011111" when X = 49 AND Y = 65 else
"110111011111" when X = 50 AND Y = 65 else
"110111011111" when X = 51 AND Y = 65 else
"110111011111" when X = 52 AND Y = 65 else
"110111011111" when X = 53 AND Y = 65 else
"110111011111" when X = 54 AND Y = 65 else
"110111011111" when X = 55 AND Y = 65 else
"110111011111" when X = 56 AND Y = 65 else
"110111011111" when X = 57 AND Y = 65 else
"110111011111" when X = 58 AND Y = 65 else
"110111011111" when X = 59 AND Y = 65 else
"110111011111" when X = 60 AND Y = 65 else
"110111011111" when X = 61 AND Y = 65 else
"110111011111" when X = 62 AND Y = 65 else
"110111011111" when X = 63 AND Y = 65 else
"110111011111" when X = 64 AND Y = 65 else
"110111011111" when X = 65 AND Y = 65 else
"110111011111" when X = 66 AND Y = 65 else
"110111011111" when X = 67 AND Y = 65 else
"110111011111" when X = 68 AND Y = 65 else
"110111011111" when X = 69 AND Y = 65 else
"110111011111" when X = 70 AND Y = 65 else
"110111011111" when X = 71 AND Y = 65 else
"110111011111" when X = 72 AND Y = 65 else
"110111011111" when X = 73 AND Y = 65 else
"110111011111" when X = 74 AND Y = 65 else
"110111011111" when X = 75 AND Y = 65 else
"110111011111" when X = 76 AND Y = 65 else
"110111011111" when X = 77 AND Y = 65 else
"110111011111" when X = 78 AND Y = 65 else
"110111011111" when X = 79 AND Y = 65 else
"110111011111" when X = 80 AND Y = 65 else
"110111011111" when X = 81 AND Y = 65 else
"110111011111" when X = 82 AND Y = 65 else
"110111011111" when X = 83 AND Y = 65 else
"110111011111" when X = 84 AND Y = 65 else
"110111011111" when X = 85 AND Y = 65 else
"110111011111" when X = 86 AND Y = 65 else
"110111011111" when X = 87 AND Y = 65 else
"110111011111" when X = 88 AND Y = 65 else
"110111011111" when X = 89 AND Y = 65 else
"110111011111" when X = 90 AND Y = 65 else
"110111011111" when X = 91 AND Y = 65 else
"110111011111" when X = 92 AND Y = 65 else
"110111011111" when X = 93 AND Y = 65 else
"110111011111" when X = 94 AND Y = 65 else
"110111011111" when X = 95 AND Y = 65 else
"110111011111" when X = 96 AND Y = 65 else
"110111011111" when X = 97 AND Y = 65 else
"110111011111" when X = 98 AND Y = 65 else
"110111011111" when X = 99 AND Y = 65 else
"110111011111" when X = 100 AND Y = 65 else
"110111011111" when X = 101 AND Y = 65 else
"110111011111" when X = 102 AND Y = 65 else
"110111011111" when X = 103 AND Y = 65 else
"110111011111" when X = 104 AND Y = 65 else
"111111111111" when X = 105 AND Y = 65 else
"111111111111" when X = 106 AND Y = 65 else
"111111111111" when X = 107 AND Y = 65 else
"111111111111" when X = 108 AND Y = 65 else
"111111111111" when X = 109 AND Y = 65 else
"111111111111" when X = 110 AND Y = 65 else
"111111111111" when X = 111 AND Y = 65 else
"111111111111" when X = 112 AND Y = 65 else
"111111111111" when X = 113 AND Y = 65 else
"111111111111" when X = 114 AND Y = 65 else
"111111111111" when X = 115 AND Y = 65 else
"111111111111" when X = 116 AND Y = 65 else
"111111111111" when X = 117 AND Y = 65 else
"111111111111" when X = 118 AND Y = 65 else
"111111111111" when X = 119 AND Y = 65 else
"111111111111" when X = 120 AND Y = 65 else
"111111111111" when X = 121 AND Y = 65 else
"111111111111" when X = 122 AND Y = 65 else
"111111111111" when X = 123 AND Y = 65 else
"111111111111" when X = 124 AND Y = 65 else
"111111111111" when X = 125 AND Y = 65 else
"111111111111" when X = 126 AND Y = 65 else
"111111111111" when X = 127 AND Y = 65 else
"111111111111" when X = 128 AND Y = 65 else
"111111111111" when X = 129 AND Y = 65 else
"111111111111" when X = 130 AND Y = 65 else
"111111111111" when X = 131 AND Y = 65 else
"111111111111" when X = 132 AND Y = 65 else
"111111111111" when X = 133 AND Y = 65 else
"111111111111" when X = 134 AND Y = 65 else
"111111111111" when X = 135 AND Y = 65 else
"111111111111" when X = 136 AND Y = 65 else
"111111111111" when X = 137 AND Y = 65 else
"111111111111" when X = 138 AND Y = 65 else
"111111111111" when X = 139 AND Y = 65 else
"111111111111" when X = 140 AND Y = 65 else
"111111111111" when X = 141 AND Y = 65 else
"111111111111" when X = 142 AND Y = 65 else
"111111111111" when X = 143 AND Y = 65 else
"111111111111" when X = 144 AND Y = 65 else
"111111111111" when X = 145 AND Y = 65 else
"111111111111" when X = 146 AND Y = 65 else
"111111111111" when X = 147 AND Y = 65 else
"111111111111" when X = 148 AND Y = 65 else
"111111111111" when X = 149 AND Y = 65 else
"111111111111" when X = 150 AND Y = 65 else
"111111111111" when X = 151 AND Y = 65 else
"111111111111" when X = 152 AND Y = 65 else
"111111111111" when X = 153 AND Y = 65 else
"111111111111" when X = 154 AND Y = 65 else
"111111111111" when X = 155 AND Y = 65 else
"111111111111" when X = 156 AND Y = 65 else
"111111111111" when X = 157 AND Y = 65 else
"111111111111" when X = 158 AND Y = 65 else
"111111111111" when X = 159 AND Y = 65 else
"111111111111" when X = 160 AND Y = 65 else
"111111111111" when X = 161 AND Y = 65 else
"111111111111" when X = 162 AND Y = 65 else
"111111111111" when X = 163 AND Y = 65 else
"111111111111" when X = 164 AND Y = 65 else
"111111111111" when X = 165 AND Y = 65 else
"111111111111" when X = 166 AND Y = 65 else
"111111111111" when X = 167 AND Y = 65 else
"111111111111" when X = 168 AND Y = 65 else
"111111111111" when X = 169 AND Y = 65 else
"111111111111" when X = 170 AND Y = 65 else
"111111111111" when X = 171 AND Y = 65 else
"111111111111" when X = 172 AND Y = 65 else
"111111111111" when X = 173 AND Y = 65 else
"111111111111" when X = 174 AND Y = 65 else
"111111111111" when X = 175 AND Y = 65 else
"111111111111" when X = 176 AND Y = 65 else
"111111111111" when X = 177 AND Y = 65 else
"111111111111" when X = 178 AND Y = 65 else
"111111111111" when X = 179 AND Y = 65 else
"111111111111" when X = 180 AND Y = 65 else
"111111111111" when X = 181 AND Y = 65 else
"111111111111" when X = 182 AND Y = 65 else
"111111111111" when X = 183 AND Y = 65 else
"111111111111" when X = 184 AND Y = 65 else
"111111111111" when X = 185 AND Y = 65 else
"111111111111" when X = 186 AND Y = 65 else
"111111111111" when X = 187 AND Y = 65 else
"111111111111" when X = 188 AND Y = 65 else
"111111111111" when X = 189 AND Y = 65 else
"111111111111" when X = 190 AND Y = 65 else
"111111111111" when X = 191 AND Y = 65 else
"111111111111" when X = 192 AND Y = 65 else
"111111111111" when X = 193 AND Y = 65 else
"111111111111" when X = 194 AND Y = 65 else
"111111111111" when X = 195 AND Y = 65 else
"111111111111" when X = 196 AND Y = 65 else
"111111111111" when X = 197 AND Y = 65 else
"111111111111" when X = 198 AND Y = 65 else
"111111111111" when X = 199 AND Y = 65 else
"111111111111" when X = 200 AND Y = 65 else
"111111111111" when X = 201 AND Y = 65 else
"111111111111" when X = 202 AND Y = 65 else
"111111111111" when X = 203 AND Y = 65 else
"111111111111" when X = 204 AND Y = 65 else
"111111111111" when X = 205 AND Y = 65 else
"111111111111" when X = 206 AND Y = 65 else
"111111111111" when X = 207 AND Y = 65 else
"111111111111" when X = 208 AND Y = 65 else
"111111111111" when X = 209 AND Y = 65 else
"111111111111" when X = 210 AND Y = 65 else
"111111111111" when X = 211 AND Y = 65 else
"111111111111" when X = 212 AND Y = 65 else
"111111111111" when X = 213 AND Y = 65 else
"111111111111" when X = 214 AND Y = 65 else
"111111111111" when X = 215 AND Y = 65 else
"111111111111" when X = 216 AND Y = 65 else
"111111111111" when X = 217 AND Y = 65 else
"111111111111" when X = 218 AND Y = 65 else
"111111111111" when X = 219 AND Y = 65 else
"111111111111" when X = 220 AND Y = 65 else
"111111111111" when X = 221 AND Y = 65 else
"111111111111" when X = 222 AND Y = 65 else
"111111111111" when X = 223 AND Y = 65 else
"111111111111" when X = 224 AND Y = 65 else
"111111111111" when X = 225 AND Y = 65 else
"111111111111" when X = 226 AND Y = 65 else
"111111111111" when X = 227 AND Y = 65 else
"111111111111" when X = 228 AND Y = 65 else
"111111111111" when X = 229 AND Y = 65 else
"111111111111" when X = 230 AND Y = 65 else
"111111111111" when X = 231 AND Y = 65 else
"111111111111" when X = 232 AND Y = 65 else
"111111111111" when X = 233 AND Y = 65 else
"111111111111" when X = 234 AND Y = 65 else
"111111111111" when X = 235 AND Y = 65 else
"111111111111" when X = 236 AND Y = 65 else
"111111111111" when X = 237 AND Y = 65 else
"111111111111" when X = 238 AND Y = 65 else
"111111111111" when X = 239 AND Y = 65 else
"111111111111" when X = 240 AND Y = 65 else
"111111111111" when X = 241 AND Y = 65 else
"111111111111" when X = 242 AND Y = 65 else
"111111111111" when X = 243 AND Y = 65 else
"111111111111" when X = 244 AND Y = 65 else
"111111111111" when X = 245 AND Y = 65 else
"111111111111" when X = 246 AND Y = 65 else
"111111111111" when X = 247 AND Y = 65 else
"111111111111" when X = 248 AND Y = 65 else
"111111111111" when X = 249 AND Y = 65 else
"111111111111" when X = 250 AND Y = 65 else
"111111111111" when X = 251 AND Y = 65 else
"111111111111" when X = 252 AND Y = 65 else
"111111111111" when X = 253 AND Y = 65 else
"111111111111" when X = 254 AND Y = 65 else
"111111111111" when X = 255 AND Y = 65 else
"111111111111" when X = 256 AND Y = 65 else
"111111111111" when X = 257 AND Y = 65 else
"111111111111" when X = 258 AND Y = 65 else
"111111111111" when X = 259 AND Y = 65 else
"111111111111" when X = 260 AND Y = 65 else
"111111111111" when X = 261 AND Y = 65 else
"111111111111" when X = 262 AND Y = 65 else
"111111111111" when X = 263 AND Y = 65 else
"111111111111" when X = 264 AND Y = 65 else
"110111011111" when X = 265 AND Y = 65 else
"110111011111" when X = 266 AND Y = 65 else
"110111011111" when X = 267 AND Y = 65 else
"110111011111" when X = 268 AND Y = 65 else
"110111011111" when X = 269 AND Y = 65 else
"110111011111" when X = 270 AND Y = 65 else
"110111011111" when X = 271 AND Y = 65 else
"110111011111" when X = 272 AND Y = 65 else
"110111011111" when X = 273 AND Y = 65 else
"110111011111" when X = 274 AND Y = 65 else
"110111011111" when X = 275 AND Y = 65 else
"110111011111" when X = 276 AND Y = 65 else
"110111011111" when X = 277 AND Y = 65 else
"110111011111" when X = 278 AND Y = 65 else
"110111011111" when X = 279 AND Y = 65 else
"000000000000" when X = 280 AND Y = 65 else
"000000000000" when X = 281 AND Y = 65 else
"000000000000" when X = 282 AND Y = 65 else
"000000000000" when X = 283 AND Y = 65 else
"000000000000" when X = 284 AND Y = 65 else
"000000000000" when X = 285 AND Y = 65 else
"000000000000" when X = 286 AND Y = 65 else
"000000000000" when X = 287 AND Y = 65 else
"000000000000" when X = 288 AND Y = 65 else
"000000000000" when X = 289 AND Y = 65 else
"000000000000" when X = 290 AND Y = 65 else
"000000000000" when X = 291 AND Y = 65 else
"000000000000" when X = 292 AND Y = 65 else
"000000000000" when X = 293 AND Y = 65 else
"000000000000" when X = 294 AND Y = 65 else
"000000000000" when X = 295 AND Y = 65 else
"000000000000" when X = 296 AND Y = 65 else
"000000000000" when X = 297 AND Y = 65 else
"000000000000" when X = 298 AND Y = 65 else
"000000000000" when X = 299 AND Y = 65 else
"000000000000" when X = 300 AND Y = 65 else
"000000000000" when X = 301 AND Y = 65 else
"000000000000" when X = 302 AND Y = 65 else
"000000000000" when X = 303 AND Y = 65 else
"000000000000" when X = 304 AND Y = 65 else
"000000000000" when X = 305 AND Y = 65 else
"000000000000" when X = 306 AND Y = 65 else
"000000000000" when X = 307 AND Y = 65 else
"000000000000" when X = 308 AND Y = 65 else
"000000000000" when X = 309 AND Y = 65 else
"000000000000" when X = 310 AND Y = 65 else
"000000000000" when X = 311 AND Y = 65 else
"000000000000" when X = 312 AND Y = 65 else
"000000000000" when X = 313 AND Y = 65 else
"000000000000" when X = 314 AND Y = 65 else
"000000000000" when X = 315 AND Y = 65 else
"000000000000" when X = 316 AND Y = 65 else
"000000000000" when X = 317 AND Y = 65 else
"000000000000" when X = 318 AND Y = 65 else
"000000000000" when X = 319 AND Y = 65 else
"000000000000" when X = 320 AND Y = 65 else
"000000000000" when X = 321 AND Y = 65 else
"000000000000" when X = 322 AND Y = 65 else
"000000000000" when X = 323 AND Y = 65 else
"000000000000" when X = 324 AND Y = 65 else
"100010011101" when X = 0 AND Y = 66 else
"100010011101" when X = 1 AND Y = 66 else
"100010011101" when X = 2 AND Y = 66 else
"100010011101" when X = 3 AND Y = 66 else
"100010011101" when X = 4 AND Y = 66 else
"100010011101" when X = 5 AND Y = 66 else
"100010011101" when X = 6 AND Y = 66 else
"100010011101" when X = 7 AND Y = 66 else
"100010011101" when X = 8 AND Y = 66 else
"100010011101" when X = 9 AND Y = 66 else
"100010011101" when X = 10 AND Y = 66 else
"100010011101" when X = 11 AND Y = 66 else
"100010011101" when X = 12 AND Y = 66 else
"100010011101" when X = 13 AND Y = 66 else
"100010011101" when X = 14 AND Y = 66 else
"100010011101" when X = 15 AND Y = 66 else
"100010011101" when X = 16 AND Y = 66 else
"100010011101" when X = 17 AND Y = 66 else
"100010011101" when X = 18 AND Y = 66 else
"100010011101" when X = 19 AND Y = 66 else
"100010011101" when X = 20 AND Y = 66 else
"100010011101" when X = 21 AND Y = 66 else
"100010011101" when X = 22 AND Y = 66 else
"100010011101" when X = 23 AND Y = 66 else
"100010011101" when X = 24 AND Y = 66 else
"100010011101" when X = 25 AND Y = 66 else
"100010011101" when X = 26 AND Y = 66 else
"100010011101" when X = 27 AND Y = 66 else
"100010011101" when X = 28 AND Y = 66 else
"100010011101" when X = 29 AND Y = 66 else
"100010011101" when X = 30 AND Y = 66 else
"100010011101" when X = 31 AND Y = 66 else
"100010011101" when X = 32 AND Y = 66 else
"100010011101" when X = 33 AND Y = 66 else
"100010011101" when X = 34 AND Y = 66 else
"110111011111" when X = 35 AND Y = 66 else
"110111011111" when X = 36 AND Y = 66 else
"110111011111" when X = 37 AND Y = 66 else
"110111011111" when X = 38 AND Y = 66 else
"110111011111" when X = 39 AND Y = 66 else
"110111011111" when X = 40 AND Y = 66 else
"110111011111" when X = 41 AND Y = 66 else
"110111011111" when X = 42 AND Y = 66 else
"110111011111" when X = 43 AND Y = 66 else
"110111011111" when X = 44 AND Y = 66 else
"110111011111" when X = 45 AND Y = 66 else
"110111011111" when X = 46 AND Y = 66 else
"110111011111" when X = 47 AND Y = 66 else
"110111011111" when X = 48 AND Y = 66 else
"110111011111" when X = 49 AND Y = 66 else
"110111011111" when X = 50 AND Y = 66 else
"110111011111" when X = 51 AND Y = 66 else
"110111011111" when X = 52 AND Y = 66 else
"110111011111" when X = 53 AND Y = 66 else
"110111011111" when X = 54 AND Y = 66 else
"110111011111" when X = 55 AND Y = 66 else
"110111011111" when X = 56 AND Y = 66 else
"110111011111" when X = 57 AND Y = 66 else
"110111011111" when X = 58 AND Y = 66 else
"110111011111" when X = 59 AND Y = 66 else
"110111011111" when X = 60 AND Y = 66 else
"110111011111" when X = 61 AND Y = 66 else
"110111011111" when X = 62 AND Y = 66 else
"110111011111" when X = 63 AND Y = 66 else
"110111011111" when X = 64 AND Y = 66 else
"110111011111" when X = 65 AND Y = 66 else
"110111011111" when X = 66 AND Y = 66 else
"110111011111" when X = 67 AND Y = 66 else
"110111011111" when X = 68 AND Y = 66 else
"110111011111" when X = 69 AND Y = 66 else
"110111011111" when X = 70 AND Y = 66 else
"110111011111" when X = 71 AND Y = 66 else
"110111011111" when X = 72 AND Y = 66 else
"110111011111" when X = 73 AND Y = 66 else
"110111011111" when X = 74 AND Y = 66 else
"110111011111" when X = 75 AND Y = 66 else
"110111011111" when X = 76 AND Y = 66 else
"110111011111" when X = 77 AND Y = 66 else
"110111011111" when X = 78 AND Y = 66 else
"110111011111" when X = 79 AND Y = 66 else
"110111011111" when X = 80 AND Y = 66 else
"110111011111" when X = 81 AND Y = 66 else
"110111011111" when X = 82 AND Y = 66 else
"110111011111" when X = 83 AND Y = 66 else
"110111011111" when X = 84 AND Y = 66 else
"110111011111" when X = 85 AND Y = 66 else
"110111011111" when X = 86 AND Y = 66 else
"110111011111" when X = 87 AND Y = 66 else
"110111011111" when X = 88 AND Y = 66 else
"110111011111" when X = 89 AND Y = 66 else
"110111011111" when X = 90 AND Y = 66 else
"110111011111" when X = 91 AND Y = 66 else
"110111011111" when X = 92 AND Y = 66 else
"110111011111" when X = 93 AND Y = 66 else
"110111011111" when X = 94 AND Y = 66 else
"110111011111" when X = 95 AND Y = 66 else
"110111011111" when X = 96 AND Y = 66 else
"110111011111" when X = 97 AND Y = 66 else
"110111011111" when X = 98 AND Y = 66 else
"110111011111" when X = 99 AND Y = 66 else
"110111011111" when X = 100 AND Y = 66 else
"110111011111" when X = 101 AND Y = 66 else
"110111011111" when X = 102 AND Y = 66 else
"110111011111" when X = 103 AND Y = 66 else
"110111011111" when X = 104 AND Y = 66 else
"111111111111" when X = 105 AND Y = 66 else
"111111111111" when X = 106 AND Y = 66 else
"111111111111" when X = 107 AND Y = 66 else
"111111111111" when X = 108 AND Y = 66 else
"111111111111" when X = 109 AND Y = 66 else
"111111111111" when X = 110 AND Y = 66 else
"111111111111" when X = 111 AND Y = 66 else
"111111111111" when X = 112 AND Y = 66 else
"111111111111" when X = 113 AND Y = 66 else
"111111111111" when X = 114 AND Y = 66 else
"111111111111" when X = 115 AND Y = 66 else
"111111111111" when X = 116 AND Y = 66 else
"111111111111" when X = 117 AND Y = 66 else
"111111111111" when X = 118 AND Y = 66 else
"111111111111" when X = 119 AND Y = 66 else
"111111111111" when X = 120 AND Y = 66 else
"111111111111" when X = 121 AND Y = 66 else
"111111111111" when X = 122 AND Y = 66 else
"111111111111" when X = 123 AND Y = 66 else
"111111111111" when X = 124 AND Y = 66 else
"111111111111" when X = 125 AND Y = 66 else
"111111111111" when X = 126 AND Y = 66 else
"111111111111" when X = 127 AND Y = 66 else
"111111111111" when X = 128 AND Y = 66 else
"111111111111" when X = 129 AND Y = 66 else
"111111111111" when X = 130 AND Y = 66 else
"111111111111" when X = 131 AND Y = 66 else
"111111111111" when X = 132 AND Y = 66 else
"111111111111" when X = 133 AND Y = 66 else
"111111111111" when X = 134 AND Y = 66 else
"111111111111" when X = 135 AND Y = 66 else
"111111111111" when X = 136 AND Y = 66 else
"111111111111" when X = 137 AND Y = 66 else
"111111111111" when X = 138 AND Y = 66 else
"111111111111" when X = 139 AND Y = 66 else
"111111111111" when X = 140 AND Y = 66 else
"111111111111" when X = 141 AND Y = 66 else
"111111111111" when X = 142 AND Y = 66 else
"111111111111" when X = 143 AND Y = 66 else
"111111111111" when X = 144 AND Y = 66 else
"111111111111" when X = 145 AND Y = 66 else
"111111111111" when X = 146 AND Y = 66 else
"111111111111" when X = 147 AND Y = 66 else
"111111111111" when X = 148 AND Y = 66 else
"111111111111" when X = 149 AND Y = 66 else
"111111111111" when X = 150 AND Y = 66 else
"111111111111" when X = 151 AND Y = 66 else
"111111111111" when X = 152 AND Y = 66 else
"111111111111" when X = 153 AND Y = 66 else
"111111111111" when X = 154 AND Y = 66 else
"111111111111" when X = 155 AND Y = 66 else
"111111111111" when X = 156 AND Y = 66 else
"111111111111" when X = 157 AND Y = 66 else
"111111111111" when X = 158 AND Y = 66 else
"111111111111" when X = 159 AND Y = 66 else
"111111111111" when X = 160 AND Y = 66 else
"111111111111" when X = 161 AND Y = 66 else
"111111111111" when X = 162 AND Y = 66 else
"111111111111" when X = 163 AND Y = 66 else
"111111111111" when X = 164 AND Y = 66 else
"111111111111" when X = 165 AND Y = 66 else
"111111111111" when X = 166 AND Y = 66 else
"111111111111" when X = 167 AND Y = 66 else
"111111111111" when X = 168 AND Y = 66 else
"111111111111" when X = 169 AND Y = 66 else
"111111111111" when X = 170 AND Y = 66 else
"111111111111" when X = 171 AND Y = 66 else
"111111111111" when X = 172 AND Y = 66 else
"111111111111" when X = 173 AND Y = 66 else
"111111111111" when X = 174 AND Y = 66 else
"111111111111" when X = 175 AND Y = 66 else
"111111111111" when X = 176 AND Y = 66 else
"111111111111" when X = 177 AND Y = 66 else
"111111111111" when X = 178 AND Y = 66 else
"111111111111" when X = 179 AND Y = 66 else
"111111111111" when X = 180 AND Y = 66 else
"111111111111" when X = 181 AND Y = 66 else
"111111111111" when X = 182 AND Y = 66 else
"111111111111" when X = 183 AND Y = 66 else
"111111111111" when X = 184 AND Y = 66 else
"111111111111" when X = 185 AND Y = 66 else
"111111111111" when X = 186 AND Y = 66 else
"111111111111" when X = 187 AND Y = 66 else
"111111111111" when X = 188 AND Y = 66 else
"111111111111" when X = 189 AND Y = 66 else
"111111111111" when X = 190 AND Y = 66 else
"111111111111" when X = 191 AND Y = 66 else
"111111111111" when X = 192 AND Y = 66 else
"111111111111" when X = 193 AND Y = 66 else
"111111111111" when X = 194 AND Y = 66 else
"111111111111" when X = 195 AND Y = 66 else
"111111111111" when X = 196 AND Y = 66 else
"111111111111" when X = 197 AND Y = 66 else
"111111111111" when X = 198 AND Y = 66 else
"111111111111" when X = 199 AND Y = 66 else
"111111111111" when X = 200 AND Y = 66 else
"111111111111" when X = 201 AND Y = 66 else
"111111111111" when X = 202 AND Y = 66 else
"111111111111" when X = 203 AND Y = 66 else
"111111111111" when X = 204 AND Y = 66 else
"111111111111" when X = 205 AND Y = 66 else
"111111111111" when X = 206 AND Y = 66 else
"111111111111" when X = 207 AND Y = 66 else
"111111111111" when X = 208 AND Y = 66 else
"111111111111" when X = 209 AND Y = 66 else
"111111111111" when X = 210 AND Y = 66 else
"111111111111" when X = 211 AND Y = 66 else
"111111111111" when X = 212 AND Y = 66 else
"111111111111" when X = 213 AND Y = 66 else
"111111111111" when X = 214 AND Y = 66 else
"111111111111" when X = 215 AND Y = 66 else
"111111111111" when X = 216 AND Y = 66 else
"111111111111" when X = 217 AND Y = 66 else
"111111111111" when X = 218 AND Y = 66 else
"111111111111" when X = 219 AND Y = 66 else
"111111111111" when X = 220 AND Y = 66 else
"111111111111" when X = 221 AND Y = 66 else
"111111111111" when X = 222 AND Y = 66 else
"111111111111" when X = 223 AND Y = 66 else
"111111111111" when X = 224 AND Y = 66 else
"111111111111" when X = 225 AND Y = 66 else
"111111111111" when X = 226 AND Y = 66 else
"111111111111" when X = 227 AND Y = 66 else
"111111111111" when X = 228 AND Y = 66 else
"111111111111" when X = 229 AND Y = 66 else
"111111111111" when X = 230 AND Y = 66 else
"111111111111" when X = 231 AND Y = 66 else
"111111111111" when X = 232 AND Y = 66 else
"111111111111" when X = 233 AND Y = 66 else
"111111111111" when X = 234 AND Y = 66 else
"111111111111" when X = 235 AND Y = 66 else
"111111111111" when X = 236 AND Y = 66 else
"111111111111" when X = 237 AND Y = 66 else
"111111111111" when X = 238 AND Y = 66 else
"111111111111" when X = 239 AND Y = 66 else
"111111111111" when X = 240 AND Y = 66 else
"111111111111" when X = 241 AND Y = 66 else
"111111111111" when X = 242 AND Y = 66 else
"111111111111" when X = 243 AND Y = 66 else
"111111111111" when X = 244 AND Y = 66 else
"111111111111" when X = 245 AND Y = 66 else
"111111111111" when X = 246 AND Y = 66 else
"111111111111" when X = 247 AND Y = 66 else
"111111111111" when X = 248 AND Y = 66 else
"111111111111" when X = 249 AND Y = 66 else
"111111111111" when X = 250 AND Y = 66 else
"111111111111" when X = 251 AND Y = 66 else
"111111111111" when X = 252 AND Y = 66 else
"111111111111" when X = 253 AND Y = 66 else
"111111111111" when X = 254 AND Y = 66 else
"111111111111" when X = 255 AND Y = 66 else
"111111111111" when X = 256 AND Y = 66 else
"111111111111" when X = 257 AND Y = 66 else
"111111111111" when X = 258 AND Y = 66 else
"111111111111" when X = 259 AND Y = 66 else
"111111111111" when X = 260 AND Y = 66 else
"111111111111" when X = 261 AND Y = 66 else
"111111111111" when X = 262 AND Y = 66 else
"111111111111" when X = 263 AND Y = 66 else
"111111111111" when X = 264 AND Y = 66 else
"110111011111" when X = 265 AND Y = 66 else
"110111011111" when X = 266 AND Y = 66 else
"110111011111" when X = 267 AND Y = 66 else
"110111011111" when X = 268 AND Y = 66 else
"110111011111" when X = 269 AND Y = 66 else
"110111011111" when X = 270 AND Y = 66 else
"110111011111" when X = 271 AND Y = 66 else
"110111011111" when X = 272 AND Y = 66 else
"110111011111" when X = 273 AND Y = 66 else
"110111011111" when X = 274 AND Y = 66 else
"110111011111" when X = 275 AND Y = 66 else
"110111011111" when X = 276 AND Y = 66 else
"110111011111" when X = 277 AND Y = 66 else
"110111011111" when X = 278 AND Y = 66 else
"110111011111" when X = 279 AND Y = 66 else
"000000000000" when X = 280 AND Y = 66 else
"000000000000" when X = 281 AND Y = 66 else
"000000000000" when X = 282 AND Y = 66 else
"000000000000" when X = 283 AND Y = 66 else
"000000000000" when X = 284 AND Y = 66 else
"000000000000" when X = 285 AND Y = 66 else
"000000000000" when X = 286 AND Y = 66 else
"000000000000" when X = 287 AND Y = 66 else
"000000000000" when X = 288 AND Y = 66 else
"000000000000" when X = 289 AND Y = 66 else
"000000000000" when X = 290 AND Y = 66 else
"000000000000" when X = 291 AND Y = 66 else
"000000000000" when X = 292 AND Y = 66 else
"000000000000" when X = 293 AND Y = 66 else
"000000000000" when X = 294 AND Y = 66 else
"000000000000" when X = 295 AND Y = 66 else
"000000000000" when X = 296 AND Y = 66 else
"000000000000" when X = 297 AND Y = 66 else
"000000000000" when X = 298 AND Y = 66 else
"000000000000" when X = 299 AND Y = 66 else
"000000000000" when X = 300 AND Y = 66 else
"000000000000" when X = 301 AND Y = 66 else
"000000000000" when X = 302 AND Y = 66 else
"000000000000" when X = 303 AND Y = 66 else
"000000000000" when X = 304 AND Y = 66 else
"000000000000" when X = 305 AND Y = 66 else
"000000000000" when X = 306 AND Y = 66 else
"000000000000" when X = 307 AND Y = 66 else
"000000000000" when X = 308 AND Y = 66 else
"000000000000" when X = 309 AND Y = 66 else
"000000000000" when X = 310 AND Y = 66 else
"000000000000" when X = 311 AND Y = 66 else
"000000000000" when X = 312 AND Y = 66 else
"000000000000" when X = 313 AND Y = 66 else
"000000000000" when X = 314 AND Y = 66 else
"000000000000" when X = 315 AND Y = 66 else
"000000000000" when X = 316 AND Y = 66 else
"000000000000" when X = 317 AND Y = 66 else
"000000000000" when X = 318 AND Y = 66 else
"000000000000" when X = 319 AND Y = 66 else
"000000000000" when X = 320 AND Y = 66 else
"000000000000" when X = 321 AND Y = 66 else
"000000000000" when X = 322 AND Y = 66 else
"000000000000" when X = 323 AND Y = 66 else
"000000000000" when X = 324 AND Y = 66 else
"100010011101" when X = 0 AND Y = 67 else
"100010011101" when X = 1 AND Y = 67 else
"100010011101" when X = 2 AND Y = 67 else
"100010011101" when X = 3 AND Y = 67 else
"100010011101" when X = 4 AND Y = 67 else
"100010011101" when X = 5 AND Y = 67 else
"100010011101" when X = 6 AND Y = 67 else
"100010011101" when X = 7 AND Y = 67 else
"100010011101" when X = 8 AND Y = 67 else
"100010011101" when X = 9 AND Y = 67 else
"100010011101" when X = 10 AND Y = 67 else
"100010011101" when X = 11 AND Y = 67 else
"100010011101" when X = 12 AND Y = 67 else
"100010011101" when X = 13 AND Y = 67 else
"100010011101" when X = 14 AND Y = 67 else
"100010011101" when X = 15 AND Y = 67 else
"100010011101" when X = 16 AND Y = 67 else
"100010011101" when X = 17 AND Y = 67 else
"100010011101" when X = 18 AND Y = 67 else
"100010011101" when X = 19 AND Y = 67 else
"100010011101" when X = 20 AND Y = 67 else
"100010011101" when X = 21 AND Y = 67 else
"100010011101" when X = 22 AND Y = 67 else
"100010011101" when X = 23 AND Y = 67 else
"100010011101" when X = 24 AND Y = 67 else
"100010011101" when X = 25 AND Y = 67 else
"100010011101" when X = 26 AND Y = 67 else
"100010011101" when X = 27 AND Y = 67 else
"100010011101" when X = 28 AND Y = 67 else
"100010011101" when X = 29 AND Y = 67 else
"100010011101" when X = 30 AND Y = 67 else
"100010011101" when X = 31 AND Y = 67 else
"100010011101" when X = 32 AND Y = 67 else
"100010011101" when X = 33 AND Y = 67 else
"100010011101" when X = 34 AND Y = 67 else
"110111011111" when X = 35 AND Y = 67 else
"110111011111" when X = 36 AND Y = 67 else
"110111011111" when X = 37 AND Y = 67 else
"110111011111" when X = 38 AND Y = 67 else
"110111011111" when X = 39 AND Y = 67 else
"110111011111" when X = 40 AND Y = 67 else
"110111011111" when X = 41 AND Y = 67 else
"110111011111" when X = 42 AND Y = 67 else
"110111011111" when X = 43 AND Y = 67 else
"110111011111" when X = 44 AND Y = 67 else
"110111011111" when X = 45 AND Y = 67 else
"110111011111" when X = 46 AND Y = 67 else
"110111011111" when X = 47 AND Y = 67 else
"110111011111" when X = 48 AND Y = 67 else
"110111011111" when X = 49 AND Y = 67 else
"110111011111" when X = 50 AND Y = 67 else
"110111011111" when X = 51 AND Y = 67 else
"110111011111" when X = 52 AND Y = 67 else
"110111011111" when X = 53 AND Y = 67 else
"110111011111" when X = 54 AND Y = 67 else
"110111011111" when X = 55 AND Y = 67 else
"110111011111" when X = 56 AND Y = 67 else
"110111011111" when X = 57 AND Y = 67 else
"110111011111" when X = 58 AND Y = 67 else
"110111011111" when X = 59 AND Y = 67 else
"110111011111" when X = 60 AND Y = 67 else
"110111011111" when X = 61 AND Y = 67 else
"110111011111" when X = 62 AND Y = 67 else
"110111011111" when X = 63 AND Y = 67 else
"110111011111" when X = 64 AND Y = 67 else
"110111011111" when X = 65 AND Y = 67 else
"110111011111" when X = 66 AND Y = 67 else
"110111011111" when X = 67 AND Y = 67 else
"110111011111" when X = 68 AND Y = 67 else
"110111011111" when X = 69 AND Y = 67 else
"110111011111" when X = 70 AND Y = 67 else
"110111011111" when X = 71 AND Y = 67 else
"110111011111" when X = 72 AND Y = 67 else
"110111011111" when X = 73 AND Y = 67 else
"110111011111" when X = 74 AND Y = 67 else
"110111011111" when X = 75 AND Y = 67 else
"110111011111" when X = 76 AND Y = 67 else
"110111011111" when X = 77 AND Y = 67 else
"110111011111" when X = 78 AND Y = 67 else
"110111011111" when X = 79 AND Y = 67 else
"110111011111" when X = 80 AND Y = 67 else
"110111011111" when X = 81 AND Y = 67 else
"110111011111" when X = 82 AND Y = 67 else
"110111011111" when X = 83 AND Y = 67 else
"110111011111" when X = 84 AND Y = 67 else
"110111011111" when X = 85 AND Y = 67 else
"110111011111" when X = 86 AND Y = 67 else
"110111011111" when X = 87 AND Y = 67 else
"110111011111" when X = 88 AND Y = 67 else
"110111011111" when X = 89 AND Y = 67 else
"110111011111" when X = 90 AND Y = 67 else
"110111011111" when X = 91 AND Y = 67 else
"110111011111" when X = 92 AND Y = 67 else
"110111011111" when X = 93 AND Y = 67 else
"110111011111" when X = 94 AND Y = 67 else
"110111011111" when X = 95 AND Y = 67 else
"110111011111" when X = 96 AND Y = 67 else
"110111011111" when X = 97 AND Y = 67 else
"110111011111" when X = 98 AND Y = 67 else
"110111011111" when X = 99 AND Y = 67 else
"110111011111" when X = 100 AND Y = 67 else
"110111011111" when X = 101 AND Y = 67 else
"110111011111" when X = 102 AND Y = 67 else
"110111011111" when X = 103 AND Y = 67 else
"110111011111" when X = 104 AND Y = 67 else
"111111111111" when X = 105 AND Y = 67 else
"111111111111" when X = 106 AND Y = 67 else
"111111111111" when X = 107 AND Y = 67 else
"111111111111" when X = 108 AND Y = 67 else
"111111111111" when X = 109 AND Y = 67 else
"111111111111" when X = 110 AND Y = 67 else
"111111111111" when X = 111 AND Y = 67 else
"111111111111" when X = 112 AND Y = 67 else
"111111111111" when X = 113 AND Y = 67 else
"111111111111" when X = 114 AND Y = 67 else
"111111111111" when X = 115 AND Y = 67 else
"111111111111" when X = 116 AND Y = 67 else
"111111111111" when X = 117 AND Y = 67 else
"111111111111" when X = 118 AND Y = 67 else
"111111111111" when X = 119 AND Y = 67 else
"111111111111" when X = 120 AND Y = 67 else
"111111111111" when X = 121 AND Y = 67 else
"111111111111" when X = 122 AND Y = 67 else
"111111111111" when X = 123 AND Y = 67 else
"111111111111" when X = 124 AND Y = 67 else
"111111111111" when X = 125 AND Y = 67 else
"111111111111" when X = 126 AND Y = 67 else
"111111111111" when X = 127 AND Y = 67 else
"111111111111" when X = 128 AND Y = 67 else
"111111111111" when X = 129 AND Y = 67 else
"111111111111" when X = 130 AND Y = 67 else
"111111111111" when X = 131 AND Y = 67 else
"111111111111" when X = 132 AND Y = 67 else
"111111111111" when X = 133 AND Y = 67 else
"111111111111" when X = 134 AND Y = 67 else
"111111111111" when X = 135 AND Y = 67 else
"111111111111" when X = 136 AND Y = 67 else
"111111111111" when X = 137 AND Y = 67 else
"111111111111" when X = 138 AND Y = 67 else
"111111111111" when X = 139 AND Y = 67 else
"111111111111" when X = 140 AND Y = 67 else
"111111111111" when X = 141 AND Y = 67 else
"111111111111" when X = 142 AND Y = 67 else
"111111111111" when X = 143 AND Y = 67 else
"111111111111" when X = 144 AND Y = 67 else
"111111111111" when X = 145 AND Y = 67 else
"111111111111" when X = 146 AND Y = 67 else
"111111111111" when X = 147 AND Y = 67 else
"111111111111" when X = 148 AND Y = 67 else
"111111111111" when X = 149 AND Y = 67 else
"111111111111" when X = 150 AND Y = 67 else
"111111111111" when X = 151 AND Y = 67 else
"111111111111" when X = 152 AND Y = 67 else
"111111111111" when X = 153 AND Y = 67 else
"111111111111" when X = 154 AND Y = 67 else
"111111111111" when X = 155 AND Y = 67 else
"111111111111" when X = 156 AND Y = 67 else
"111111111111" when X = 157 AND Y = 67 else
"111111111111" when X = 158 AND Y = 67 else
"111111111111" when X = 159 AND Y = 67 else
"111111111111" when X = 160 AND Y = 67 else
"111111111111" when X = 161 AND Y = 67 else
"111111111111" when X = 162 AND Y = 67 else
"111111111111" when X = 163 AND Y = 67 else
"111111111111" when X = 164 AND Y = 67 else
"111111111111" when X = 165 AND Y = 67 else
"111111111111" when X = 166 AND Y = 67 else
"111111111111" when X = 167 AND Y = 67 else
"111111111111" when X = 168 AND Y = 67 else
"111111111111" when X = 169 AND Y = 67 else
"111111111111" when X = 170 AND Y = 67 else
"111111111111" when X = 171 AND Y = 67 else
"111111111111" when X = 172 AND Y = 67 else
"111111111111" when X = 173 AND Y = 67 else
"111111111111" when X = 174 AND Y = 67 else
"111111111111" when X = 175 AND Y = 67 else
"111111111111" when X = 176 AND Y = 67 else
"111111111111" when X = 177 AND Y = 67 else
"111111111111" when X = 178 AND Y = 67 else
"111111111111" when X = 179 AND Y = 67 else
"111111111111" when X = 180 AND Y = 67 else
"111111111111" when X = 181 AND Y = 67 else
"111111111111" when X = 182 AND Y = 67 else
"111111111111" when X = 183 AND Y = 67 else
"111111111111" when X = 184 AND Y = 67 else
"111111111111" when X = 185 AND Y = 67 else
"111111111111" when X = 186 AND Y = 67 else
"111111111111" when X = 187 AND Y = 67 else
"111111111111" when X = 188 AND Y = 67 else
"111111111111" when X = 189 AND Y = 67 else
"111111111111" when X = 190 AND Y = 67 else
"111111111111" when X = 191 AND Y = 67 else
"111111111111" when X = 192 AND Y = 67 else
"111111111111" when X = 193 AND Y = 67 else
"111111111111" when X = 194 AND Y = 67 else
"111111111111" when X = 195 AND Y = 67 else
"111111111111" when X = 196 AND Y = 67 else
"111111111111" when X = 197 AND Y = 67 else
"111111111111" when X = 198 AND Y = 67 else
"111111111111" when X = 199 AND Y = 67 else
"111111111111" when X = 200 AND Y = 67 else
"111111111111" when X = 201 AND Y = 67 else
"111111111111" when X = 202 AND Y = 67 else
"111111111111" when X = 203 AND Y = 67 else
"111111111111" when X = 204 AND Y = 67 else
"111111111111" when X = 205 AND Y = 67 else
"111111111111" when X = 206 AND Y = 67 else
"111111111111" when X = 207 AND Y = 67 else
"111111111111" when X = 208 AND Y = 67 else
"111111111111" when X = 209 AND Y = 67 else
"111111111111" when X = 210 AND Y = 67 else
"111111111111" when X = 211 AND Y = 67 else
"111111111111" when X = 212 AND Y = 67 else
"111111111111" when X = 213 AND Y = 67 else
"111111111111" when X = 214 AND Y = 67 else
"111111111111" when X = 215 AND Y = 67 else
"111111111111" when X = 216 AND Y = 67 else
"111111111111" when X = 217 AND Y = 67 else
"111111111111" when X = 218 AND Y = 67 else
"111111111111" when X = 219 AND Y = 67 else
"111111111111" when X = 220 AND Y = 67 else
"111111111111" when X = 221 AND Y = 67 else
"111111111111" when X = 222 AND Y = 67 else
"111111111111" when X = 223 AND Y = 67 else
"111111111111" when X = 224 AND Y = 67 else
"111111111111" when X = 225 AND Y = 67 else
"111111111111" when X = 226 AND Y = 67 else
"111111111111" when X = 227 AND Y = 67 else
"111111111111" when X = 228 AND Y = 67 else
"111111111111" when X = 229 AND Y = 67 else
"111111111111" when X = 230 AND Y = 67 else
"111111111111" when X = 231 AND Y = 67 else
"111111111111" when X = 232 AND Y = 67 else
"111111111111" when X = 233 AND Y = 67 else
"111111111111" when X = 234 AND Y = 67 else
"111111111111" when X = 235 AND Y = 67 else
"111111111111" when X = 236 AND Y = 67 else
"111111111111" when X = 237 AND Y = 67 else
"111111111111" when X = 238 AND Y = 67 else
"111111111111" when X = 239 AND Y = 67 else
"111111111111" when X = 240 AND Y = 67 else
"111111111111" when X = 241 AND Y = 67 else
"111111111111" when X = 242 AND Y = 67 else
"111111111111" when X = 243 AND Y = 67 else
"111111111111" when X = 244 AND Y = 67 else
"111111111111" when X = 245 AND Y = 67 else
"111111111111" when X = 246 AND Y = 67 else
"111111111111" when X = 247 AND Y = 67 else
"111111111111" when X = 248 AND Y = 67 else
"111111111111" when X = 249 AND Y = 67 else
"111111111111" when X = 250 AND Y = 67 else
"111111111111" when X = 251 AND Y = 67 else
"111111111111" when X = 252 AND Y = 67 else
"111111111111" when X = 253 AND Y = 67 else
"111111111111" when X = 254 AND Y = 67 else
"111111111111" when X = 255 AND Y = 67 else
"111111111111" when X = 256 AND Y = 67 else
"111111111111" when X = 257 AND Y = 67 else
"111111111111" when X = 258 AND Y = 67 else
"111111111111" when X = 259 AND Y = 67 else
"111111111111" when X = 260 AND Y = 67 else
"111111111111" when X = 261 AND Y = 67 else
"111111111111" when X = 262 AND Y = 67 else
"111111111111" when X = 263 AND Y = 67 else
"111111111111" when X = 264 AND Y = 67 else
"110111011111" when X = 265 AND Y = 67 else
"110111011111" when X = 266 AND Y = 67 else
"110111011111" when X = 267 AND Y = 67 else
"110111011111" when X = 268 AND Y = 67 else
"110111011111" when X = 269 AND Y = 67 else
"110111011111" when X = 270 AND Y = 67 else
"110111011111" when X = 271 AND Y = 67 else
"110111011111" when X = 272 AND Y = 67 else
"110111011111" when X = 273 AND Y = 67 else
"110111011111" when X = 274 AND Y = 67 else
"110111011111" when X = 275 AND Y = 67 else
"110111011111" when X = 276 AND Y = 67 else
"110111011111" when X = 277 AND Y = 67 else
"110111011111" when X = 278 AND Y = 67 else
"110111011111" when X = 279 AND Y = 67 else
"000000000000" when X = 280 AND Y = 67 else
"000000000000" when X = 281 AND Y = 67 else
"000000000000" when X = 282 AND Y = 67 else
"000000000000" when X = 283 AND Y = 67 else
"000000000000" when X = 284 AND Y = 67 else
"000000000000" when X = 285 AND Y = 67 else
"000000000000" when X = 286 AND Y = 67 else
"000000000000" when X = 287 AND Y = 67 else
"000000000000" when X = 288 AND Y = 67 else
"000000000000" when X = 289 AND Y = 67 else
"000000000000" when X = 290 AND Y = 67 else
"000000000000" when X = 291 AND Y = 67 else
"000000000000" when X = 292 AND Y = 67 else
"000000000000" when X = 293 AND Y = 67 else
"000000000000" when X = 294 AND Y = 67 else
"000000000000" when X = 295 AND Y = 67 else
"000000000000" when X = 296 AND Y = 67 else
"000000000000" when X = 297 AND Y = 67 else
"000000000000" when X = 298 AND Y = 67 else
"000000000000" when X = 299 AND Y = 67 else
"000000000000" when X = 300 AND Y = 67 else
"000000000000" when X = 301 AND Y = 67 else
"000000000000" when X = 302 AND Y = 67 else
"000000000000" when X = 303 AND Y = 67 else
"000000000000" when X = 304 AND Y = 67 else
"000000000000" when X = 305 AND Y = 67 else
"000000000000" when X = 306 AND Y = 67 else
"000000000000" when X = 307 AND Y = 67 else
"000000000000" when X = 308 AND Y = 67 else
"000000000000" when X = 309 AND Y = 67 else
"000000000000" when X = 310 AND Y = 67 else
"000000000000" when X = 311 AND Y = 67 else
"000000000000" when X = 312 AND Y = 67 else
"000000000000" when X = 313 AND Y = 67 else
"000000000000" when X = 314 AND Y = 67 else
"000000000000" when X = 315 AND Y = 67 else
"000000000000" when X = 316 AND Y = 67 else
"000000000000" when X = 317 AND Y = 67 else
"000000000000" when X = 318 AND Y = 67 else
"000000000000" when X = 319 AND Y = 67 else
"000000000000" when X = 320 AND Y = 67 else
"000000000000" when X = 321 AND Y = 67 else
"000000000000" when X = 322 AND Y = 67 else
"000000000000" when X = 323 AND Y = 67 else
"000000000000" when X = 324 AND Y = 67 else
"100010011101" when X = 0 AND Y = 68 else
"100010011101" when X = 1 AND Y = 68 else
"100010011101" when X = 2 AND Y = 68 else
"100010011101" when X = 3 AND Y = 68 else
"100010011101" when X = 4 AND Y = 68 else
"100010011101" when X = 5 AND Y = 68 else
"100010011101" when X = 6 AND Y = 68 else
"100010011101" when X = 7 AND Y = 68 else
"100010011101" when X = 8 AND Y = 68 else
"100010011101" when X = 9 AND Y = 68 else
"100010011101" when X = 10 AND Y = 68 else
"100010011101" when X = 11 AND Y = 68 else
"100010011101" when X = 12 AND Y = 68 else
"100010011101" when X = 13 AND Y = 68 else
"100010011101" when X = 14 AND Y = 68 else
"100010011101" when X = 15 AND Y = 68 else
"100010011101" when X = 16 AND Y = 68 else
"100010011101" when X = 17 AND Y = 68 else
"100010011101" when X = 18 AND Y = 68 else
"100010011101" when X = 19 AND Y = 68 else
"100010011101" when X = 20 AND Y = 68 else
"100010011101" when X = 21 AND Y = 68 else
"100010011101" when X = 22 AND Y = 68 else
"100010011101" when X = 23 AND Y = 68 else
"100010011101" when X = 24 AND Y = 68 else
"100010011101" when X = 25 AND Y = 68 else
"100010011101" when X = 26 AND Y = 68 else
"100010011101" when X = 27 AND Y = 68 else
"100010011101" when X = 28 AND Y = 68 else
"100010011101" when X = 29 AND Y = 68 else
"100010011101" when X = 30 AND Y = 68 else
"100010011101" when X = 31 AND Y = 68 else
"100010011101" when X = 32 AND Y = 68 else
"100010011101" when X = 33 AND Y = 68 else
"100010011101" when X = 34 AND Y = 68 else
"110111011111" when X = 35 AND Y = 68 else
"110111011111" when X = 36 AND Y = 68 else
"110111011111" when X = 37 AND Y = 68 else
"110111011111" when X = 38 AND Y = 68 else
"110111011111" when X = 39 AND Y = 68 else
"110111011111" when X = 40 AND Y = 68 else
"110111011111" when X = 41 AND Y = 68 else
"110111011111" when X = 42 AND Y = 68 else
"110111011111" when X = 43 AND Y = 68 else
"110111011111" when X = 44 AND Y = 68 else
"110111011111" when X = 45 AND Y = 68 else
"110111011111" when X = 46 AND Y = 68 else
"110111011111" when X = 47 AND Y = 68 else
"110111011111" when X = 48 AND Y = 68 else
"110111011111" when X = 49 AND Y = 68 else
"110111011111" when X = 50 AND Y = 68 else
"110111011111" when X = 51 AND Y = 68 else
"110111011111" when X = 52 AND Y = 68 else
"110111011111" when X = 53 AND Y = 68 else
"110111011111" when X = 54 AND Y = 68 else
"110111011111" when X = 55 AND Y = 68 else
"110111011111" when X = 56 AND Y = 68 else
"110111011111" when X = 57 AND Y = 68 else
"110111011111" when X = 58 AND Y = 68 else
"110111011111" when X = 59 AND Y = 68 else
"110111011111" when X = 60 AND Y = 68 else
"110111011111" when X = 61 AND Y = 68 else
"110111011111" when X = 62 AND Y = 68 else
"110111011111" when X = 63 AND Y = 68 else
"110111011111" when X = 64 AND Y = 68 else
"110111011111" when X = 65 AND Y = 68 else
"110111011111" when X = 66 AND Y = 68 else
"110111011111" when X = 67 AND Y = 68 else
"110111011111" when X = 68 AND Y = 68 else
"110111011111" when X = 69 AND Y = 68 else
"110111011111" when X = 70 AND Y = 68 else
"110111011111" when X = 71 AND Y = 68 else
"110111011111" when X = 72 AND Y = 68 else
"110111011111" when X = 73 AND Y = 68 else
"110111011111" when X = 74 AND Y = 68 else
"110111011111" when X = 75 AND Y = 68 else
"110111011111" when X = 76 AND Y = 68 else
"110111011111" when X = 77 AND Y = 68 else
"110111011111" when X = 78 AND Y = 68 else
"110111011111" when X = 79 AND Y = 68 else
"110111011111" when X = 80 AND Y = 68 else
"110111011111" when X = 81 AND Y = 68 else
"110111011111" when X = 82 AND Y = 68 else
"110111011111" when X = 83 AND Y = 68 else
"110111011111" when X = 84 AND Y = 68 else
"110111011111" when X = 85 AND Y = 68 else
"110111011111" when X = 86 AND Y = 68 else
"110111011111" when X = 87 AND Y = 68 else
"110111011111" when X = 88 AND Y = 68 else
"110111011111" when X = 89 AND Y = 68 else
"110111011111" when X = 90 AND Y = 68 else
"110111011111" when X = 91 AND Y = 68 else
"110111011111" when X = 92 AND Y = 68 else
"110111011111" when X = 93 AND Y = 68 else
"110111011111" when X = 94 AND Y = 68 else
"110111011111" when X = 95 AND Y = 68 else
"110111011111" when X = 96 AND Y = 68 else
"110111011111" when X = 97 AND Y = 68 else
"110111011111" when X = 98 AND Y = 68 else
"110111011111" when X = 99 AND Y = 68 else
"110111011111" when X = 100 AND Y = 68 else
"110111011111" when X = 101 AND Y = 68 else
"110111011111" when X = 102 AND Y = 68 else
"110111011111" when X = 103 AND Y = 68 else
"110111011111" when X = 104 AND Y = 68 else
"111111111111" when X = 105 AND Y = 68 else
"111111111111" when X = 106 AND Y = 68 else
"111111111111" when X = 107 AND Y = 68 else
"111111111111" when X = 108 AND Y = 68 else
"111111111111" when X = 109 AND Y = 68 else
"111111111111" when X = 110 AND Y = 68 else
"111111111111" when X = 111 AND Y = 68 else
"111111111111" when X = 112 AND Y = 68 else
"111111111111" when X = 113 AND Y = 68 else
"111111111111" when X = 114 AND Y = 68 else
"111111111111" when X = 115 AND Y = 68 else
"111111111111" when X = 116 AND Y = 68 else
"111111111111" when X = 117 AND Y = 68 else
"111111111111" when X = 118 AND Y = 68 else
"111111111111" when X = 119 AND Y = 68 else
"111111111111" when X = 120 AND Y = 68 else
"111111111111" when X = 121 AND Y = 68 else
"111111111111" when X = 122 AND Y = 68 else
"111111111111" when X = 123 AND Y = 68 else
"111111111111" when X = 124 AND Y = 68 else
"111111111111" when X = 125 AND Y = 68 else
"111111111111" when X = 126 AND Y = 68 else
"111111111111" when X = 127 AND Y = 68 else
"111111111111" when X = 128 AND Y = 68 else
"111111111111" when X = 129 AND Y = 68 else
"111111111111" when X = 130 AND Y = 68 else
"111111111111" when X = 131 AND Y = 68 else
"111111111111" when X = 132 AND Y = 68 else
"111111111111" when X = 133 AND Y = 68 else
"111111111111" when X = 134 AND Y = 68 else
"111111111111" when X = 135 AND Y = 68 else
"111111111111" when X = 136 AND Y = 68 else
"111111111111" when X = 137 AND Y = 68 else
"111111111111" when X = 138 AND Y = 68 else
"111111111111" when X = 139 AND Y = 68 else
"111111111111" when X = 140 AND Y = 68 else
"111111111111" when X = 141 AND Y = 68 else
"111111111111" when X = 142 AND Y = 68 else
"111111111111" when X = 143 AND Y = 68 else
"111111111111" when X = 144 AND Y = 68 else
"111111111111" when X = 145 AND Y = 68 else
"111111111111" when X = 146 AND Y = 68 else
"111111111111" when X = 147 AND Y = 68 else
"111111111111" when X = 148 AND Y = 68 else
"111111111111" when X = 149 AND Y = 68 else
"111111111111" when X = 150 AND Y = 68 else
"111111111111" when X = 151 AND Y = 68 else
"111111111111" when X = 152 AND Y = 68 else
"111111111111" when X = 153 AND Y = 68 else
"111111111111" when X = 154 AND Y = 68 else
"111111111111" when X = 155 AND Y = 68 else
"111111111111" when X = 156 AND Y = 68 else
"111111111111" when X = 157 AND Y = 68 else
"111111111111" when X = 158 AND Y = 68 else
"111111111111" when X = 159 AND Y = 68 else
"111111111111" when X = 160 AND Y = 68 else
"111111111111" when X = 161 AND Y = 68 else
"111111111111" when X = 162 AND Y = 68 else
"111111111111" when X = 163 AND Y = 68 else
"111111111111" when X = 164 AND Y = 68 else
"111111111111" when X = 165 AND Y = 68 else
"111111111111" when X = 166 AND Y = 68 else
"111111111111" when X = 167 AND Y = 68 else
"111111111111" when X = 168 AND Y = 68 else
"111111111111" when X = 169 AND Y = 68 else
"111111111111" when X = 170 AND Y = 68 else
"111111111111" when X = 171 AND Y = 68 else
"111111111111" when X = 172 AND Y = 68 else
"111111111111" when X = 173 AND Y = 68 else
"111111111111" when X = 174 AND Y = 68 else
"111111111111" when X = 175 AND Y = 68 else
"111111111111" when X = 176 AND Y = 68 else
"111111111111" when X = 177 AND Y = 68 else
"111111111111" when X = 178 AND Y = 68 else
"111111111111" when X = 179 AND Y = 68 else
"111111111111" when X = 180 AND Y = 68 else
"111111111111" when X = 181 AND Y = 68 else
"111111111111" when X = 182 AND Y = 68 else
"111111111111" when X = 183 AND Y = 68 else
"111111111111" when X = 184 AND Y = 68 else
"111111111111" when X = 185 AND Y = 68 else
"111111111111" when X = 186 AND Y = 68 else
"111111111111" when X = 187 AND Y = 68 else
"111111111111" when X = 188 AND Y = 68 else
"111111111111" when X = 189 AND Y = 68 else
"111111111111" when X = 190 AND Y = 68 else
"111111111111" when X = 191 AND Y = 68 else
"111111111111" when X = 192 AND Y = 68 else
"111111111111" when X = 193 AND Y = 68 else
"111111111111" when X = 194 AND Y = 68 else
"111111111111" when X = 195 AND Y = 68 else
"111111111111" when X = 196 AND Y = 68 else
"111111111111" when X = 197 AND Y = 68 else
"111111111111" when X = 198 AND Y = 68 else
"111111111111" when X = 199 AND Y = 68 else
"111111111111" when X = 200 AND Y = 68 else
"111111111111" when X = 201 AND Y = 68 else
"111111111111" when X = 202 AND Y = 68 else
"111111111111" when X = 203 AND Y = 68 else
"111111111111" when X = 204 AND Y = 68 else
"111111111111" when X = 205 AND Y = 68 else
"111111111111" when X = 206 AND Y = 68 else
"111111111111" when X = 207 AND Y = 68 else
"111111111111" when X = 208 AND Y = 68 else
"111111111111" when X = 209 AND Y = 68 else
"111111111111" when X = 210 AND Y = 68 else
"111111111111" when X = 211 AND Y = 68 else
"111111111111" when X = 212 AND Y = 68 else
"111111111111" when X = 213 AND Y = 68 else
"111111111111" when X = 214 AND Y = 68 else
"111111111111" when X = 215 AND Y = 68 else
"111111111111" when X = 216 AND Y = 68 else
"111111111111" when X = 217 AND Y = 68 else
"111111111111" when X = 218 AND Y = 68 else
"111111111111" when X = 219 AND Y = 68 else
"111111111111" when X = 220 AND Y = 68 else
"111111111111" when X = 221 AND Y = 68 else
"111111111111" when X = 222 AND Y = 68 else
"111111111111" when X = 223 AND Y = 68 else
"111111111111" when X = 224 AND Y = 68 else
"111111111111" when X = 225 AND Y = 68 else
"111111111111" when X = 226 AND Y = 68 else
"111111111111" when X = 227 AND Y = 68 else
"111111111111" when X = 228 AND Y = 68 else
"111111111111" when X = 229 AND Y = 68 else
"111111111111" when X = 230 AND Y = 68 else
"111111111111" when X = 231 AND Y = 68 else
"111111111111" when X = 232 AND Y = 68 else
"111111111111" when X = 233 AND Y = 68 else
"111111111111" when X = 234 AND Y = 68 else
"111111111111" when X = 235 AND Y = 68 else
"111111111111" when X = 236 AND Y = 68 else
"111111111111" when X = 237 AND Y = 68 else
"111111111111" when X = 238 AND Y = 68 else
"111111111111" when X = 239 AND Y = 68 else
"111111111111" when X = 240 AND Y = 68 else
"111111111111" when X = 241 AND Y = 68 else
"111111111111" when X = 242 AND Y = 68 else
"111111111111" when X = 243 AND Y = 68 else
"111111111111" when X = 244 AND Y = 68 else
"111111111111" when X = 245 AND Y = 68 else
"111111111111" when X = 246 AND Y = 68 else
"111111111111" when X = 247 AND Y = 68 else
"111111111111" when X = 248 AND Y = 68 else
"111111111111" when X = 249 AND Y = 68 else
"111111111111" when X = 250 AND Y = 68 else
"111111111111" when X = 251 AND Y = 68 else
"111111111111" when X = 252 AND Y = 68 else
"111111111111" when X = 253 AND Y = 68 else
"111111111111" when X = 254 AND Y = 68 else
"111111111111" when X = 255 AND Y = 68 else
"111111111111" when X = 256 AND Y = 68 else
"111111111111" when X = 257 AND Y = 68 else
"111111111111" when X = 258 AND Y = 68 else
"111111111111" when X = 259 AND Y = 68 else
"111111111111" when X = 260 AND Y = 68 else
"111111111111" when X = 261 AND Y = 68 else
"111111111111" when X = 262 AND Y = 68 else
"111111111111" when X = 263 AND Y = 68 else
"111111111111" when X = 264 AND Y = 68 else
"110111011111" when X = 265 AND Y = 68 else
"110111011111" when X = 266 AND Y = 68 else
"110111011111" when X = 267 AND Y = 68 else
"110111011111" when X = 268 AND Y = 68 else
"110111011111" when X = 269 AND Y = 68 else
"110111011111" when X = 270 AND Y = 68 else
"110111011111" when X = 271 AND Y = 68 else
"110111011111" when X = 272 AND Y = 68 else
"110111011111" when X = 273 AND Y = 68 else
"110111011111" when X = 274 AND Y = 68 else
"110111011111" when X = 275 AND Y = 68 else
"110111011111" when X = 276 AND Y = 68 else
"110111011111" when X = 277 AND Y = 68 else
"110111011111" when X = 278 AND Y = 68 else
"110111011111" when X = 279 AND Y = 68 else
"000000000000" when X = 280 AND Y = 68 else
"000000000000" when X = 281 AND Y = 68 else
"000000000000" when X = 282 AND Y = 68 else
"000000000000" when X = 283 AND Y = 68 else
"000000000000" when X = 284 AND Y = 68 else
"000000000000" when X = 285 AND Y = 68 else
"000000000000" when X = 286 AND Y = 68 else
"000000000000" when X = 287 AND Y = 68 else
"000000000000" when X = 288 AND Y = 68 else
"000000000000" when X = 289 AND Y = 68 else
"000000000000" when X = 290 AND Y = 68 else
"000000000000" when X = 291 AND Y = 68 else
"000000000000" when X = 292 AND Y = 68 else
"000000000000" when X = 293 AND Y = 68 else
"000000000000" when X = 294 AND Y = 68 else
"000000000000" when X = 295 AND Y = 68 else
"000000000000" when X = 296 AND Y = 68 else
"000000000000" when X = 297 AND Y = 68 else
"000000000000" when X = 298 AND Y = 68 else
"000000000000" when X = 299 AND Y = 68 else
"000000000000" when X = 300 AND Y = 68 else
"000000000000" when X = 301 AND Y = 68 else
"000000000000" when X = 302 AND Y = 68 else
"000000000000" when X = 303 AND Y = 68 else
"000000000000" when X = 304 AND Y = 68 else
"000000000000" when X = 305 AND Y = 68 else
"000000000000" when X = 306 AND Y = 68 else
"000000000000" when X = 307 AND Y = 68 else
"000000000000" when X = 308 AND Y = 68 else
"000000000000" when X = 309 AND Y = 68 else
"000000000000" when X = 310 AND Y = 68 else
"000000000000" when X = 311 AND Y = 68 else
"000000000000" when X = 312 AND Y = 68 else
"000000000000" when X = 313 AND Y = 68 else
"000000000000" when X = 314 AND Y = 68 else
"000000000000" when X = 315 AND Y = 68 else
"000000000000" when X = 316 AND Y = 68 else
"000000000000" when X = 317 AND Y = 68 else
"000000000000" when X = 318 AND Y = 68 else
"000000000000" when X = 319 AND Y = 68 else
"000000000000" when X = 320 AND Y = 68 else
"000000000000" when X = 321 AND Y = 68 else
"000000000000" when X = 322 AND Y = 68 else
"000000000000" when X = 323 AND Y = 68 else
"000000000000" when X = 324 AND Y = 68 else
"100010011101" when X = 0 AND Y = 69 else
"100010011101" when X = 1 AND Y = 69 else
"100010011101" when X = 2 AND Y = 69 else
"100010011101" when X = 3 AND Y = 69 else
"100010011101" when X = 4 AND Y = 69 else
"100010011101" when X = 5 AND Y = 69 else
"100010011101" when X = 6 AND Y = 69 else
"100010011101" when X = 7 AND Y = 69 else
"100010011101" when X = 8 AND Y = 69 else
"100010011101" when X = 9 AND Y = 69 else
"100010011101" when X = 10 AND Y = 69 else
"100010011101" when X = 11 AND Y = 69 else
"100010011101" when X = 12 AND Y = 69 else
"100010011101" when X = 13 AND Y = 69 else
"100010011101" when X = 14 AND Y = 69 else
"100010011101" when X = 15 AND Y = 69 else
"100010011101" when X = 16 AND Y = 69 else
"100010011101" when X = 17 AND Y = 69 else
"100010011101" when X = 18 AND Y = 69 else
"100010011101" when X = 19 AND Y = 69 else
"100010011101" when X = 20 AND Y = 69 else
"100010011101" when X = 21 AND Y = 69 else
"100010011101" when X = 22 AND Y = 69 else
"100010011101" when X = 23 AND Y = 69 else
"100010011101" when X = 24 AND Y = 69 else
"100010011101" when X = 25 AND Y = 69 else
"100010011101" when X = 26 AND Y = 69 else
"100010011101" when X = 27 AND Y = 69 else
"100010011101" when X = 28 AND Y = 69 else
"100010011101" when X = 29 AND Y = 69 else
"100010011101" when X = 30 AND Y = 69 else
"100010011101" when X = 31 AND Y = 69 else
"100010011101" when X = 32 AND Y = 69 else
"100010011101" when X = 33 AND Y = 69 else
"100010011101" when X = 34 AND Y = 69 else
"110111011111" when X = 35 AND Y = 69 else
"110111011111" when X = 36 AND Y = 69 else
"110111011111" when X = 37 AND Y = 69 else
"110111011111" when X = 38 AND Y = 69 else
"110111011111" when X = 39 AND Y = 69 else
"110111011111" when X = 40 AND Y = 69 else
"110111011111" when X = 41 AND Y = 69 else
"110111011111" when X = 42 AND Y = 69 else
"110111011111" when X = 43 AND Y = 69 else
"110111011111" when X = 44 AND Y = 69 else
"110111011111" when X = 45 AND Y = 69 else
"110111011111" when X = 46 AND Y = 69 else
"110111011111" when X = 47 AND Y = 69 else
"110111011111" when X = 48 AND Y = 69 else
"110111011111" when X = 49 AND Y = 69 else
"110111011111" when X = 50 AND Y = 69 else
"110111011111" when X = 51 AND Y = 69 else
"110111011111" when X = 52 AND Y = 69 else
"110111011111" when X = 53 AND Y = 69 else
"110111011111" when X = 54 AND Y = 69 else
"110111011111" when X = 55 AND Y = 69 else
"110111011111" when X = 56 AND Y = 69 else
"110111011111" when X = 57 AND Y = 69 else
"110111011111" when X = 58 AND Y = 69 else
"110111011111" when X = 59 AND Y = 69 else
"110111011111" when X = 60 AND Y = 69 else
"110111011111" when X = 61 AND Y = 69 else
"110111011111" when X = 62 AND Y = 69 else
"110111011111" when X = 63 AND Y = 69 else
"110111011111" when X = 64 AND Y = 69 else
"110111011111" when X = 65 AND Y = 69 else
"110111011111" when X = 66 AND Y = 69 else
"110111011111" when X = 67 AND Y = 69 else
"110111011111" when X = 68 AND Y = 69 else
"110111011111" when X = 69 AND Y = 69 else
"110111011111" when X = 70 AND Y = 69 else
"110111011111" when X = 71 AND Y = 69 else
"110111011111" when X = 72 AND Y = 69 else
"110111011111" when X = 73 AND Y = 69 else
"110111011111" when X = 74 AND Y = 69 else
"110111011111" when X = 75 AND Y = 69 else
"110111011111" when X = 76 AND Y = 69 else
"110111011111" when X = 77 AND Y = 69 else
"110111011111" when X = 78 AND Y = 69 else
"110111011111" when X = 79 AND Y = 69 else
"110111011111" when X = 80 AND Y = 69 else
"110111011111" when X = 81 AND Y = 69 else
"110111011111" when X = 82 AND Y = 69 else
"110111011111" when X = 83 AND Y = 69 else
"110111011111" when X = 84 AND Y = 69 else
"110111011111" when X = 85 AND Y = 69 else
"110111011111" when X = 86 AND Y = 69 else
"110111011111" when X = 87 AND Y = 69 else
"110111011111" when X = 88 AND Y = 69 else
"110111011111" when X = 89 AND Y = 69 else
"110111011111" when X = 90 AND Y = 69 else
"110111011111" when X = 91 AND Y = 69 else
"110111011111" when X = 92 AND Y = 69 else
"110111011111" when X = 93 AND Y = 69 else
"110111011111" when X = 94 AND Y = 69 else
"110111011111" when X = 95 AND Y = 69 else
"110111011111" when X = 96 AND Y = 69 else
"110111011111" when X = 97 AND Y = 69 else
"110111011111" when X = 98 AND Y = 69 else
"110111011111" when X = 99 AND Y = 69 else
"110111011111" when X = 100 AND Y = 69 else
"110111011111" when X = 101 AND Y = 69 else
"110111011111" when X = 102 AND Y = 69 else
"110111011111" when X = 103 AND Y = 69 else
"110111011111" when X = 104 AND Y = 69 else
"111111111111" when X = 105 AND Y = 69 else
"111111111111" when X = 106 AND Y = 69 else
"111111111111" when X = 107 AND Y = 69 else
"111111111111" when X = 108 AND Y = 69 else
"111111111111" when X = 109 AND Y = 69 else
"111111111111" when X = 110 AND Y = 69 else
"111111111111" when X = 111 AND Y = 69 else
"111111111111" when X = 112 AND Y = 69 else
"111111111111" when X = 113 AND Y = 69 else
"111111111111" when X = 114 AND Y = 69 else
"111111111111" when X = 115 AND Y = 69 else
"111111111111" when X = 116 AND Y = 69 else
"111111111111" when X = 117 AND Y = 69 else
"111111111111" when X = 118 AND Y = 69 else
"111111111111" when X = 119 AND Y = 69 else
"111111111111" when X = 120 AND Y = 69 else
"111111111111" when X = 121 AND Y = 69 else
"111111111111" when X = 122 AND Y = 69 else
"111111111111" when X = 123 AND Y = 69 else
"111111111111" when X = 124 AND Y = 69 else
"111111111111" when X = 125 AND Y = 69 else
"111111111111" when X = 126 AND Y = 69 else
"111111111111" when X = 127 AND Y = 69 else
"111111111111" when X = 128 AND Y = 69 else
"111111111111" when X = 129 AND Y = 69 else
"111111111111" when X = 130 AND Y = 69 else
"111111111111" when X = 131 AND Y = 69 else
"111111111111" when X = 132 AND Y = 69 else
"111111111111" when X = 133 AND Y = 69 else
"111111111111" when X = 134 AND Y = 69 else
"111111111111" when X = 135 AND Y = 69 else
"111111111111" when X = 136 AND Y = 69 else
"111111111111" when X = 137 AND Y = 69 else
"111111111111" when X = 138 AND Y = 69 else
"111111111111" when X = 139 AND Y = 69 else
"111111111111" when X = 140 AND Y = 69 else
"111111111111" when X = 141 AND Y = 69 else
"111111111111" when X = 142 AND Y = 69 else
"111111111111" when X = 143 AND Y = 69 else
"111111111111" when X = 144 AND Y = 69 else
"111111111111" when X = 145 AND Y = 69 else
"111111111111" when X = 146 AND Y = 69 else
"111111111111" when X = 147 AND Y = 69 else
"111111111111" when X = 148 AND Y = 69 else
"111111111111" when X = 149 AND Y = 69 else
"111111111111" when X = 150 AND Y = 69 else
"111111111111" when X = 151 AND Y = 69 else
"111111111111" when X = 152 AND Y = 69 else
"111111111111" when X = 153 AND Y = 69 else
"111111111111" when X = 154 AND Y = 69 else
"111111111111" when X = 155 AND Y = 69 else
"111111111111" when X = 156 AND Y = 69 else
"111111111111" when X = 157 AND Y = 69 else
"111111111111" when X = 158 AND Y = 69 else
"111111111111" when X = 159 AND Y = 69 else
"111111111111" when X = 160 AND Y = 69 else
"111111111111" when X = 161 AND Y = 69 else
"111111111111" when X = 162 AND Y = 69 else
"111111111111" when X = 163 AND Y = 69 else
"111111111111" when X = 164 AND Y = 69 else
"111111111111" when X = 165 AND Y = 69 else
"111111111111" when X = 166 AND Y = 69 else
"111111111111" when X = 167 AND Y = 69 else
"111111111111" when X = 168 AND Y = 69 else
"111111111111" when X = 169 AND Y = 69 else
"111111111111" when X = 170 AND Y = 69 else
"111111111111" when X = 171 AND Y = 69 else
"111111111111" when X = 172 AND Y = 69 else
"111111111111" when X = 173 AND Y = 69 else
"111111111111" when X = 174 AND Y = 69 else
"111111111111" when X = 175 AND Y = 69 else
"111111111111" when X = 176 AND Y = 69 else
"111111111111" when X = 177 AND Y = 69 else
"111111111111" when X = 178 AND Y = 69 else
"111111111111" when X = 179 AND Y = 69 else
"111111111111" when X = 180 AND Y = 69 else
"111111111111" when X = 181 AND Y = 69 else
"111111111111" when X = 182 AND Y = 69 else
"111111111111" when X = 183 AND Y = 69 else
"111111111111" when X = 184 AND Y = 69 else
"111111111111" when X = 185 AND Y = 69 else
"111111111111" when X = 186 AND Y = 69 else
"111111111111" when X = 187 AND Y = 69 else
"111111111111" when X = 188 AND Y = 69 else
"111111111111" when X = 189 AND Y = 69 else
"111111111111" when X = 190 AND Y = 69 else
"111111111111" when X = 191 AND Y = 69 else
"111111111111" when X = 192 AND Y = 69 else
"111111111111" when X = 193 AND Y = 69 else
"111111111111" when X = 194 AND Y = 69 else
"111111111111" when X = 195 AND Y = 69 else
"111111111111" when X = 196 AND Y = 69 else
"111111111111" when X = 197 AND Y = 69 else
"111111111111" when X = 198 AND Y = 69 else
"111111111111" when X = 199 AND Y = 69 else
"111111111111" when X = 200 AND Y = 69 else
"111111111111" when X = 201 AND Y = 69 else
"111111111111" when X = 202 AND Y = 69 else
"111111111111" when X = 203 AND Y = 69 else
"111111111111" when X = 204 AND Y = 69 else
"111111111111" when X = 205 AND Y = 69 else
"111111111111" when X = 206 AND Y = 69 else
"111111111111" when X = 207 AND Y = 69 else
"111111111111" when X = 208 AND Y = 69 else
"111111111111" when X = 209 AND Y = 69 else
"111111111111" when X = 210 AND Y = 69 else
"111111111111" when X = 211 AND Y = 69 else
"111111111111" when X = 212 AND Y = 69 else
"111111111111" when X = 213 AND Y = 69 else
"111111111111" when X = 214 AND Y = 69 else
"111111111111" when X = 215 AND Y = 69 else
"111111111111" when X = 216 AND Y = 69 else
"111111111111" when X = 217 AND Y = 69 else
"111111111111" when X = 218 AND Y = 69 else
"111111111111" when X = 219 AND Y = 69 else
"111111111111" when X = 220 AND Y = 69 else
"111111111111" when X = 221 AND Y = 69 else
"111111111111" when X = 222 AND Y = 69 else
"111111111111" when X = 223 AND Y = 69 else
"111111111111" when X = 224 AND Y = 69 else
"111111111111" when X = 225 AND Y = 69 else
"111111111111" when X = 226 AND Y = 69 else
"111111111111" when X = 227 AND Y = 69 else
"111111111111" when X = 228 AND Y = 69 else
"111111111111" when X = 229 AND Y = 69 else
"111111111111" when X = 230 AND Y = 69 else
"111111111111" when X = 231 AND Y = 69 else
"111111111111" when X = 232 AND Y = 69 else
"111111111111" when X = 233 AND Y = 69 else
"111111111111" when X = 234 AND Y = 69 else
"111111111111" when X = 235 AND Y = 69 else
"111111111111" when X = 236 AND Y = 69 else
"111111111111" when X = 237 AND Y = 69 else
"111111111111" when X = 238 AND Y = 69 else
"111111111111" when X = 239 AND Y = 69 else
"111111111111" when X = 240 AND Y = 69 else
"111111111111" when X = 241 AND Y = 69 else
"111111111111" when X = 242 AND Y = 69 else
"111111111111" when X = 243 AND Y = 69 else
"111111111111" when X = 244 AND Y = 69 else
"111111111111" when X = 245 AND Y = 69 else
"111111111111" when X = 246 AND Y = 69 else
"111111111111" when X = 247 AND Y = 69 else
"111111111111" when X = 248 AND Y = 69 else
"111111111111" when X = 249 AND Y = 69 else
"111111111111" when X = 250 AND Y = 69 else
"111111111111" when X = 251 AND Y = 69 else
"111111111111" when X = 252 AND Y = 69 else
"111111111111" when X = 253 AND Y = 69 else
"111111111111" when X = 254 AND Y = 69 else
"111111111111" when X = 255 AND Y = 69 else
"111111111111" when X = 256 AND Y = 69 else
"111111111111" when X = 257 AND Y = 69 else
"111111111111" when X = 258 AND Y = 69 else
"111111111111" when X = 259 AND Y = 69 else
"111111111111" when X = 260 AND Y = 69 else
"111111111111" when X = 261 AND Y = 69 else
"111111111111" when X = 262 AND Y = 69 else
"111111111111" when X = 263 AND Y = 69 else
"111111111111" when X = 264 AND Y = 69 else
"110111011111" when X = 265 AND Y = 69 else
"110111011111" when X = 266 AND Y = 69 else
"110111011111" when X = 267 AND Y = 69 else
"110111011111" when X = 268 AND Y = 69 else
"110111011111" when X = 269 AND Y = 69 else
"110111011111" when X = 270 AND Y = 69 else
"110111011111" when X = 271 AND Y = 69 else
"110111011111" when X = 272 AND Y = 69 else
"110111011111" when X = 273 AND Y = 69 else
"110111011111" when X = 274 AND Y = 69 else
"110111011111" when X = 275 AND Y = 69 else
"110111011111" when X = 276 AND Y = 69 else
"110111011111" when X = 277 AND Y = 69 else
"110111011111" when X = 278 AND Y = 69 else
"110111011111" when X = 279 AND Y = 69 else
"000000000000" when X = 280 AND Y = 69 else
"000000000000" when X = 281 AND Y = 69 else
"000000000000" when X = 282 AND Y = 69 else
"000000000000" when X = 283 AND Y = 69 else
"000000000000" when X = 284 AND Y = 69 else
"000000000000" when X = 285 AND Y = 69 else
"000000000000" when X = 286 AND Y = 69 else
"000000000000" when X = 287 AND Y = 69 else
"000000000000" when X = 288 AND Y = 69 else
"000000000000" when X = 289 AND Y = 69 else
"000000000000" when X = 290 AND Y = 69 else
"000000000000" when X = 291 AND Y = 69 else
"000000000000" when X = 292 AND Y = 69 else
"000000000000" when X = 293 AND Y = 69 else
"000000000000" when X = 294 AND Y = 69 else
"000000000000" when X = 295 AND Y = 69 else
"000000000000" when X = 296 AND Y = 69 else
"000000000000" when X = 297 AND Y = 69 else
"000000000000" when X = 298 AND Y = 69 else
"000000000000" when X = 299 AND Y = 69 else
"000000000000" when X = 300 AND Y = 69 else
"000000000000" when X = 301 AND Y = 69 else
"000000000000" when X = 302 AND Y = 69 else
"000000000000" when X = 303 AND Y = 69 else
"000000000000" when X = 304 AND Y = 69 else
"000000000000" when X = 305 AND Y = 69 else
"000000000000" when X = 306 AND Y = 69 else
"000000000000" when X = 307 AND Y = 69 else
"000000000000" when X = 308 AND Y = 69 else
"000000000000" when X = 309 AND Y = 69 else
"000000000000" when X = 310 AND Y = 69 else
"000000000000" when X = 311 AND Y = 69 else
"000000000000" when X = 312 AND Y = 69 else
"000000000000" when X = 313 AND Y = 69 else
"000000000000" when X = 314 AND Y = 69 else
"000000000000" when X = 315 AND Y = 69 else
"000000000000" when X = 316 AND Y = 69 else
"000000000000" when X = 317 AND Y = 69 else
"000000000000" when X = 318 AND Y = 69 else
"000000000000" when X = 319 AND Y = 69 else
"000000000000" when X = 320 AND Y = 69 else
"000000000000" when X = 321 AND Y = 69 else
"000000000000" when X = 322 AND Y = 69 else
"000000000000" when X = 323 AND Y = 69 else
"000000000000" when X = 324 AND Y = 69 else
"100010011101" when X = 0 AND Y = 70 else
"100010011101" when X = 1 AND Y = 70 else
"100010011101" when X = 2 AND Y = 70 else
"100010011101" when X = 3 AND Y = 70 else
"100010011101" when X = 4 AND Y = 70 else
"100010011101" when X = 5 AND Y = 70 else
"100010011101" when X = 6 AND Y = 70 else
"100010011101" when X = 7 AND Y = 70 else
"100010011101" when X = 8 AND Y = 70 else
"100010011101" when X = 9 AND Y = 70 else
"100010011101" when X = 10 AND Y = 70 else
"100010011101" when X = 11 AND Y = 70 else
"100010011101" when X = 12 AND Y = 70 else
"100010011101" when X = 13 AND Y = 70 else
"100010011101" when X = 14 AND Y = 70 else
"100010011101" when X = 15 AND Y = 70 else
"100010011101" when X = 16 AND Y = 70 else
"100010011101" when X = 17 AND Y = 70 else
"100010011101" when X = 18 AND Y = 70 else
"100010011101" when X = 19 AND Y = 70 else
"100010011101" when X = 20 AND Y = 70 else
"100010011101" when X = 21 AND Y = 70 else
"100010011101" when X = 22 AND Y = 70 else
"100010011101" when X = 23 AND Y = 70 else
"100010011101" when X = 24 AND Y = 70 else
"100010011101" when X = 25 AND Y = 70 else
"100010011101" when X = 26 AND Y = 70 else
"100010011101" when X = 27 AND Y = 70 else
"100010011101" when X = 28 AND Y = 70 else
"100010011101" when X = 29 AND Y = 70 else
"110111011111" when X = 30 AND Y = 70 else
"110111011111" when X = 31 AND Y = 70 else
"110111011111" when X = 32 AND Y = 70 else
"110111011111" when X = 33 AND Y = 70 else
"110111011111" when X = 34 AND Y = 70 else
"110111011111" when X = 35 AND Y = 70 else
"110111011111" when X = 36 AND Y = 70 else
"110111011111" when X = 37 AND Y = 70 else
"110111011111" when X = 38 AND Y = 70 else
"110111011111" when X = 39 AND Y = 70 else
"110111011111" when X = 40 AND Y = 70 else
"110111011111" when X = 41 AND Y = 70 else
"110111011111" when X = 42 AND Y = 70 else
"110111011111" when X = 43 AND Y = 70 else
"110111011111" when X = 44 AND Y = 70 else
"110111011111" when X = 45 AND Y = 70 else
"110111011111" when X = 46 AND Y = 70 else
"110111011111" when X = 47 AND Y = 70 else
"110111011111" when X = 48 AND Y = 70 else
"110111011111" when X = 49 AND Y = 70 else
"110111011111" when X = 50 AND Y = 70 else
"110111011111" when X = 51 AND Y = 70 else
"110111011111" when X = 52 AND Y = 70 else
"110111011111" when X = 53 AND Y = 70 else
"110111011111" when X = 54 AND Y = 70 else
"110111011111" when X = 55 AND Y = 70 else
"110111011111" when X = 56 AND Y = 70 else
"110111011111" when X = 57 AND Y = 70 else
"110111011111" when X = 58 AND Y = 70 else
"110111011111" when X = 59 AND Y = 70 else
"110111011111" when X = 60 AND Y = 70 else
"110111011111" when X = 61 AND Y = 70 else
"110111011111" when X = 62 AND Y = 70 else
"110111011111" when X = 63 AND Y = 70 else
"110111011111" when X = 64 AND Y = 70 else
"110111011111" when X = 65 AND Y = 70 else
"110111011111" when X = 66 AND Y = 70 else
"110111011111" when X = 67 AND Y = 70 else
"110111011111" when X = 68 AND Y = 70 else
"110111011111" when X = 69 AND Y = 70 else
"110111011111" when X = 70 AND Y = 70 else
"110111011111" when X = 71 AND Y = 70 else
"110111011111" when X = 72 AND Y = 70 else
"110111011111" when X = 73 AND Y = 70 else
"110111011111" when X = 74 AND Y = 70 else
"110111011111" when X = 75 AND Y = 70 else
"110111011111" when X = 76 AND Y = 70 else
"110111011111" when X = 77 AND Y = 70 else
"110111011111" when X = 78 AND Y = 70 else
"110111011111" when X = 79 AND Y = 70 else
"110111011111" when X = 80 AND Y = 70 else
"110111011111" when X = 81 AND Y = 70 else
"110111011111" when X = 82 AND Y = 70 else
"110111011111" when X = 83 AND Y = 70 else
"110111011111" when X = 84 AND Y = 70 else
"110111011111" when X = 85 AND Y = 70 else
"110111011111" when X = 86 AND Y = 70 else
"110111011111" when X = 87 AND Y = 70 else
"110111011111" when X = 88 AND Y = 70 else
"110111011111" when X = 89 AND Y = 70 else
"110111011111" when X = 90 AND Y = 70 else
"110111011111" when X = 91 AND Y = 70 else
"110111011111" when X = 92 AND Y = 70 else
"110111011111" when X = 93 AND Y = 70 else
"110111011111" when X = 94 AND Y = 70 else
"110111011111" when X = 95 AND Y = 70 else
"110111011111" when X = 96 AND Y = 70 else
"110111011111" when X = 97 AND Y = 70 else
"110111011111" when X = 98 AND Y = 70 else
"110111011111" when X = 99 AND Y = 70 else
"110111011111" when X = 100 AND Y = 70 else
"110111011111" when X = 101 AND Y = 70 else
"110111011111" when X = 102 AND Y = 70 else
"110111011111" when X = 103 AND Y = 70 else
"110111011111" when X = 104 AND Y = 70 else
"111111111111" when X = 105 AND Y = 70 else
"111111111111" when X = 106 AND Y = 70 else
"111111111111" when X = 107 AND Y = 70 else
"111111111111" when X = 108 AND Y = 70 else
"111111111111" when X = 109 AND Y = 70 else
"111111111111" when X = 110 AND Y = 70 else
"111111111111" when X = 111 AND Y = 70 else
"111111111111" when X = 112 AND Y = 70 else
"111111111111" when X = 113 AND Y = 70 else
"111111111111" when X = 114 AND Y = 70 else
"111111111111" when X = 115 AND Y = 70 else
"111111111111" when X = 116 AND Y = 70 else
"111111111111" when X = 117 AND Y = 70 else
"111111111111" when X = 118 AND Y = 70 else
"111111111111" when X = 119 AND Y = 70 else
"111111111111" when X = 120 AND Y = 70 else
"111111111111" when X = 121 AND Y = 70 else
"111111111111" when X = 122 AND Y = 70 else
"111111111111" when X = 123 AND Y = 70 else
"111111111111" when X = 124 AND Y = 70 else
"111111111111" when X = 125 AND Y = 70 else
"111111111111" when X = 126 AND Y = 70 else
"111111111111" when X = 127 AND Y = 70 else
"111111111111" when X = 128 AND Y = 70 else
"111111111111" when X = 129 AND Y = 70 else
"111111111111" when X = 130 AND Y = 70 else
"111111111111" when X = 131 AND Y = 70 else
"111111111111" when X = 132 AND Y = 70 else
"111111111111" when X = 133 AND Y = 70 else
"111111111111" when X = 134 AND Y = 70 else
"111111111111" when X = 135 AND Y = 70 else
"111111111111" when X = 136 AND Y = 70 else
"111111111111" when X = 137 AND Y = 70 else
"111111111111" when X = 138 AND Y = 70 else
"111111111111" when X = 139 AND Y = 70 else
"111111111111" when X = 140 AND Y = 70 else
"111111111111" when X = 141 AND Y = 70 else
"111111111111" when X = 142 AND Y = 70 else
"111111111111" when X = 143 AND Y = 70 else
"111111111111" when X = 144 AND Y = 70 else
"111111111111" when X = 145 AND Y = 70 else
"111111111111" when X = 146 AND Y = 70 else
"111111111111" when X = 147 AND Y = 70 else
"111111111111" when X = 148 AND Y = 70 else
"111111111111" when X = 149 AND Y = 70 else
"111111111111" when X = 150 AND Y = 70 else
"111111111111" when X = 151 AND Y = 70 else
"111111111111" when X = 152 AND Y = 70 else
"111111111111" when X = 153 AND Y = 70 else
"111111111111" when X = 154 AND Y = 70 else
"111111111111" when X = 155 AND Y = 70 else
"111111111111" when X = 156 AND Y = 70 else
"111111111111" when X = 157 AND Y = 70 else
"111111111111" when X = 158 AND Y = 70 else
"111111111111" when X = 159 AND Y = 70 else
"111111111111" when X = 160 AND Y = 70 else
"111111111111" when X = 161 AND Y = 70 else
"111111111111" when X = 162 AND Y = 70 else
"111111111111" when X = 163 AND Y = 70 else
"111111111111" when X = 164 AND Y = 70 else
"111111111111" when X = 165 AND Y = 70 else
"111111111111" when X = 166 AND Y = 70 else
"111111111111" when X = 167 AND Y = 70 else
"111111111111" when X = 168 AND Y = 70 else
"111111111111" when X = 169 AND Y = 70 else
"111111111111" when X = 170 AND Y = 70 else
"111111111111" when X = 171 AND Y = 70 else
"111111111111" when X = 172 AND Y = 70 else
"111111111111" when X = 173 AND Y = 70 else
"111111111111" when X = 174 AND Y = 70 else
"111111111111" when X = 175 AND Y = 70 else
"111111111111" when X = 176 AND Y = 70 else
"111111111111" when X = 177 AND Y = 70 else
"111111111111" when X = 178 AND Y = 70 else
"111111111111" when X = 179 AND Y = 70 else
"111111111111" when X = 180 AND Y = 70 else
"111111111111" when X = 181 AND Y = 70 else
"111111111111" when X = 182 AND Y = 70 else
"111111111111" when X = 183 AND Y = 70 else
"111111111111" when X = 184 AND Y = 70 else
"111111111111" when X = 185 AND Y = 70 else
"111111111111" when X = 186 AND Y = 70 else
"111111111111" when X = 187 AND Y = 70 else
"111111111111" when X = 188 AND Y = 70 else
"111111111111" when X = 189 AND Y = 70 else
"111111111111" when X = 190 AND Y = 70 else
"111111111111" when X = 191 AND Y = 70 else
"111111111111" when X = 192 AND Y = 70 else
"111111111111" when X = 193 AND Y = 70 else
"111111111111" when X = 194 AND Y = 70 else
"111111111111" when X = 195 AND Y = 70 else
"111111111111" when X = 196 AND Y = 70 else
"111111111111" when X = 197 AND Y = 70 else
"111111111111" when X = 198 AND Y = 70 else
"111111111111" when X = 199 AND Y = 70 else
"111111111111" when X = 200 AND Y = 70 else
"111111111111" when X = 201 AND Y = 70 else
"111111111111" when X = 202 AND Y = 70 else
"111111111111" when X = 203 AND Y = 70 else
"111111111111" when X = 204 AND Y = 70 else
"111111111111" when X = 205 AND Y = 70 else
"111111111111" when X = 206 AND Y = 70 else
"111111111111" when X = 207 AND Y = 70 else
"111111111111" when X = 208 AND Y = 70 else
"111111111111" when X = 209 AND Y = 70 else
"111111111111" when X = 210 AND Y = 70 else
"111111111111" when X = 211 AND Y = 70 else
"111111111111" when X = 212 AND Y = 70 else
"111111111111" when X = 213 AND Y = 70 else
"111111111111" when X = 214 AND Y = 70 else
"111111111111" when X = 215 AND Y = 70 else
"111111111111" when X = 216 AND Y = 70 else
"111111111111" when X = 217 AND Y = 70 else
"111111111111" when X = 218 AND Y = 70 else
"111111111111" when X = 219 AND Y = 70 else
"111111111111" when X = 220 AND Y = 70 else
"111111111111" when X = 221 AND Y = 70 else
"111111111111" when X = 222 AND Y = 70 else
"111111111111" when X = 223 AND Y = 70 else
"111111111111" when X = 224 AND Y = 70 else
"111111111111" when X = 225 AND Y = 70 else
"111111111111" when X = 226 AND Y = 70 else
"111111111111" when X = 227 AND Y = 70 else
"111111111111" when X = 228 AND Y = 70 else
"111111111111" when X = 229 AND Y = 70 else
"111111111111" when X = 230 AND Y = 70 else
"111111111111" when X = 231 AND Y = 70 else
"111111111111" when X = 232 AND Y = 70 else
"111111111111" when X = 233 AND Y = 70 else
"111111111111" when X = 234 AND Y = 70 else
"111111111111" when X = 235 AND Y = 70 else
"111111111111" when X = 236 AND Y = 70 else
"111111111111" when X = 237 AND Y = 70 else
"111111111111" when X = 238 AND Y = 70 else
"111111111111" when X = 239 AND Y = 70 else
"111111111111" when X = 240 AND Y = 70 else
"111111111111" when X = 241 AND Y = 70 else
"111111111111" when X = 242 AND Y = 70 else
"111111111111" when X = 243 AND Y = 70 else
"111111111111" when X = 244 AND Y = 70 else
"111111111111" when X = 245 AND Y = 70 else
"111111111111" when X = 246 AND Y = 70 else
"111111111111" when X = 247 AND Y = 70 else
"111111111111" when X = 248 AND Y = 70 else
"111111111111" when X = 249 AND Y = 70 else
"111111111111" when X = 250 AND Y = 70 else
"111111111111" when X = 251 AND Y = 70 else
"111111111111" when X = 252 AND Y = 70 else
"111111111111" when X = 253 AND Y = 70 else
"111111111111" when X = 254 AND Y = 70 else
"111111111111" when X = 255 AND Y = 70 else
"111111111111" when X = 256 AND Y = 70 else
"111111111111" when X = 257 AND Y = 70 else
"111111111111" when X = 258 AND Y = 70 else
"111111111111" when X = 259 AND Y = 70 else
"111111111111" when X = 260 AND Y = 70 else
"111111111111" when X = 261 AND Y = 70 else
"111111111111" when X = 262 AND Y = 70 else
"111111111111" when X = 263 AND Y = 70 else
"111111111111" when X = 264 AND Y = 70 else
"110111011111" when X = 265 AND Y = 70 else
"110111011111" when X = 266 AND Y = 70 else
"110111011111" when X = 267 AND Y = 70 else
"110111011111" when X = 268 AND Y = 70 else
"110111011111" when X = 269 AND Y = 70 else
"110111011111" when X = 270 AND Y = 70 else
"110111011111" when X = 271 AND Y = 70 else
"110111011111" when X = 272 AND Y = 70 else
"110111011111" when X = 273 AND Y = 70 else
"110111011111" when X = 274 AND Y = 70 else
"110111011111" when X = 275 AND Y = 70 else
"110111011111" when X = 276 AND Y = 70 else
"110111011111" when X = 277 AND Y = 70 else
"110111011111" when X = 278 AND Y = 70 else
"110111011111" when X = 279 AND Y = 70 else
"000000000000" when X = 280 AND Y = 70 else
"000000000000" when X = 281 AND Y = 70 else
"000000000000" when X = 282 AND Y = 70 else
"000000000000" when X = 283 AND Y = 70 else
"000000000000" when X = 284 AND Y = 70 else
"000000000000" when X = 285 AND Y = 70 else
"000000000000" when X = 286 AND Y = 70 else
"000000000000" when X = 287 AND Y = 70 else
"000000000000" when X = 288 AND Y = 70 else
"000000000000" when X = 289 AND Y = 70 else
"000000000000" when X = 290 AND Y = 70 else
"000000000000" when X = 291 AND Y = 70 else
"000000000000" when X = 292 AND Y = 70 else
"000000000000" when X = 293 AND Y = 70 else
"000000000000" when X = 294 AND Y = 70 else
"000000000000" when X = 295 AND Y = 70 else
"000000000000" when X = 296 AND Y = 70 else
"000000000000" when X = 297 AND Y = 70 else
"000000000000" when X = 298 AND Y = 70 else
"000000000000" when X = 299 AND Y = 70 else
"000000000000" when X = 300 AND Y = 70 else
"000000000000" when X = 301 AND Y = 70 else
"000000000000" when X = 302 AND Y = 70 else
"000000000000" when X = 303 AND Y = 70 else
"000000000000" when X = 304 AND Y = 70 else
"000000000000" when X = 305 AND Y = 70 else
"000000000000" when X = 306 AND Y = 70 else
"000000000000" when X = 307 AND Y = 70 else
"000000000000" when X = 308 AND Y = 70 else
"000000000000" when X = 309 AND Y = 70 else
"000000000000" when X = 310 AND Y = 70 else
"000000000000" when X = 311 AND Y = 70 else
"000000000000" when X = 312 AND Y = 70 else
"000000000000" when X = 313 AND Y = 70 else
"000000000000" when X = 314 AND Y = 70 else
"000000000000" when X = 315 AND Y = 70 else
"000000000000" when X = 316 AND Y = 70 else
"000000000000" when X = 317 AND Y = 70 else
"000000000000" when X = 318 AND Y = 70 else
"000000000000" when X = 319 AND Y = 70 else
"000000000000" when X = 320 AND Y = 70 else
"000000000000" when X = 321 AND Y = 70 else
"000000000000" when X = 322 AND Y = 70 else
"000000000000" when X = 323 AND Y = 70 else
"000000000000" when X = 324 AND Y = 70 else
"100010011101" when X = 0 AND Y = 71 else
"100010011101" when X = 1 AND Y = 71 else
"100010011101" when X = 2 AND Y = 71 else
"100010011101" when X = 3 AND Y = 71 else
"100010011101" when X = 4 AND Y = 71 else
"100010011101" when X = 5 AND Y = 71 else
"100010011101" when X = 6 AND Y = 71 else
"100010011101" when X = 7 AND Y = 71 else
"100010011101" when X = 8 AND Y = 71 else
"100010011101" when X = 9 AND Y = 71 else
"100010011101" when X = 10 AND Y = 71 else
"100010011101" when X = 11 AND Y = 71 else
"100010011101" when X = 12 AND Y = 71 else
"100010011101" when X = 13 AND Y = 71 else
"100010011101" when X = 14 AND Y = 71 else
"100010011101" when X = 15 AND Y = 71 else
"100010011101" when X = 16 AND Y = 71 else
"100010011101" when X = 17 AND Y = 71 else
"100010011101" when X = 18 AND Y = 71 else
"100010011101" when X = 19 AND Y = 71 else
"100010011101" when X = 20 AND Y = 71 else
"100010011101" when X = 21 AND Y = 71 else
"100010011101" when X = 22 AND Y = 71 else
"100010011101" when X = 23 AND Y = 71 else
"100010011101" when X = 24 AND Y = 71 else
"100010011101" when X = 25 AND Y = 71 else
"100010011101" when X = 26 AND Y = 71 else
"100010011101" when X = 27 AND Y = 71 else
"100010011101" when X = 28 AND Y = 71 else
"100010011101" when X = 29 AND Y = 71 else
"110111011111" when X = 30 AND Y = 71 else
"110111011111" when X = 31 AND Y = 71 else
"110111011111" when X = 32 AND Y = 71 else
"110111011111" when X = 33 AND Y = 71 else
"110111011111" when X = 34 AND Y = 71 else
"110111011111" when X = 35 AND Y = 71 else
"110111011111" when X = 36 AND Y = 71 else
"110111011111" when X = 37 AND Y = 71 else
"110111011111" when X = 38 AND Y = 71 else
"110111011111" when X = 39 AND Y = 71 else
"110111011111" when X = 40 AND Y = 71 else
"110111011111" when X = 41 AND Y = 71 else
"110111011111" when X = 42 AND Y = 71 else
"110111011111" when X = 43 AND Y = 71 else
"110111011111" when X = 44 AND Y = 71 else
"110111011111" when X = 45 AND Y = 71 else
"110111011111" when X = 46 AND Y = 71 else
"110111011111" when X = 47 AND Y = 71 else
"110111011111" when X = 48 AND Y = 71 else
"110111011111" when X = 49 AND Y = 71 else
"110111011111" when X = 50 AND Y = 71 else
"110111011111" when X = 51 AND Y = 71 else
"110111011111" when X = 52 AND Y = 71 else
"110111011111" when X = 53 AND Y = 71 else
"110111011111" when X = 54 AND Y = 71 else
"110111011111" when X = 55 AND Y = 71 else
"110111011111" when X = 56 AND Y = 71 else
"110111011111" when X = 57 AND Y = 71 else
"110111011111" when X = 58 AND Y = 71 else
"110111011111" when X = 59 AND Y = 71 else
"110111011111" when X = 60 AND Y = 71 else
"110111011111" when X = 61 AND Y = 71 else
"110111011111" when X = 62 AND Y = 71 else
"110111011111" when X = 63 AND Y = 71 else
"110111011111" when X = 64 AND Y = 71 else
"110111011111" when X = 65 AND Y = 71 else
"110111011111" when X = 66 AND Y = 71 else
"110111011111" when X = 67 AND Y = 71 else
"110111011111" when X = 68 AND Y = 71 else
"110111011111" when X = 69 AND Y = 71 else
"110111011111" when X = 70 AND Y = 71 else
"110111011111" when X = 71 AND Y = 71 else
"110111011111" when X = 72 AND Y = 71 else
"110111011111" when X = 73 AND Y = 71 else
"110111011111" when X = 74 AND Y = 71 else
"110111011111" when X = 75 AND Y = 71 else
"110111011111" when X = 76 AND Y = 71 else
"110111011111" when X = 77 AND Y = 71 else
"110111011111" when X = 78 AND Y = 71 else
"110111011111" when X = 79 AND Y = 71 else
"110111011111" when X = 80 AND Y = 71 else
"110111011111" when X = 81 AND Y = 71 else
"110111011111" when X = 82 AND Y = 71 else
"110111011111" when X = 83 AND Y = 71 else
"110111011111" when X = 84 AND Y = 71 else
"110111011111" when X = 85 AND Y = 71 else
"110111011111" when X = 86 AND Y = 71 else
"110111011111" when X = 87 AND Y = 71 else
"110111011111" when X = 88 AND Y = 71 else
"110111011111" when X = 89 AND Y = 71 else
"110111011111" when X = 90 AND Y = 71 else
"110111011111" when X = 91 AND Y = 71 else
"110111011111" when X = 92 AND Y = 71 else
"110111011111" when X = 93 AND Y = 71 else
"110111011111" when X = 94 AND Y = 71 else
"110111011111" when X = 95 AND Y = 71 else
"110111011111" when X = 96 AND Y = 71 else
"110111011111" when X = 97 AND Y = 71 else
"110111011111" when X = 98 AND Y = 71 else
"110111011111" when X = 99 AND Y = 71 else
"110111011111" when X = 100 AND Y = 71 else
"110111011111" when X = 101 AND Y = 71 else
"110111011111" when X = 102 AND Y = 71 else
"110111011111" when X = 103 AND Y = 71 else
"110111011111" when X = 104 AND Y = 71 else
"111111111111" when X = 105 AND Y = 71 else
"111111111111" when X = 106 AND Y = 71 else
"111111111111" when X = 107 AND Y = 71 else
"111111111111" when X = 108 AND Y = 71 else
"111111111111" when X = 109 AND Y = 71 else
"111111111111" when X = 110 AND Y = 71 else
"111111111111" when X = 111 AND Y = 71 else
"111111111111" when X = 112 AND Y = 71 else
"111111111111" when X = 113 AND Y = 71 else
"111111111111" when X = 114 AND Y = 71 else
"111111111111" when X = 115 AND Y = 71 else
"111111111111" when X = 116 AND Y = 71 else
"111111111111" when X = 117 AND Y = 71 else
"111111111111" when X = 118 AND Y = 71 else
"111111111111" when X = 119 AND Y = 71 else
"111111111111" when X = 120 AND Y = 71 else
"111111111111" when X = 121 AND Y = 71 else
"111111111111" when X = 122 AND Y = 71 else
"111111111111" when X = 123 AND Y = 71 else
"111111111111" when X = 124 AND Y = 71 else
"111111111111" when X = 125 AND Y = 71 else
"111111111111" when X = 126 AND Y = 71 else
"111111111111" when X = 127 AND Y = 71 else
"111111111111" when X = 128 AND Y = 71 else
"111111111111" when X = 129 AND Y = 71 else
"111111111111" when X = 130 AND Y = 71 else
"111111111111" when X = 131 AND Y = 71 else
"111111111111" when X = 132 AND Y = 71 else
"111111111111" when X = 133 AND Y = 71 else
"111111111111" when X = 134 AND Y = 71 else
"111111111111" when X = 135 AND Y = 71 else
"111111111111" when X = 136 AND Y = 71 else
"111111111111" when X = 137 AND Y = 71 else
"111111111111" when X = 138 AND Y = 71 else
"111111111111" when X = 139 AND Y = 71 else
"111111111111" when X = 140 AND Y = 71 else
"111111111111" when X = 141 AND Y = 71 else
"111111111111" when X = 142 AND Y = 71 else
"111111111111" when X = 143 AND Y = 71 else
"111111111111" when X = 144 AND Y = 71 else
"111111111111" when X = 145 AND Y = 71 else
"111111111111" when X = 146 AND Y = 71 else
"111111111111" when X = 147 AND Y = 71 else
"111111111111" when X = 148 AND Y = 71 else
"111111111111" when X = 149 AND Y = 71 else
"111111111111" when X = 150 AND Y = 71 else
"111111111111" when X = 151 AND Y = 71 else
"111111111111" when X = 152 AND Y = 71 else
"111111111111" when X = 153 AND Y = 71 else
"111111111111" when X = 154 AND Y = 71 else
"111111111111" when X = 155 AND Y = 71 else
"111111111111" when X = 156 AND Y = 71 else
"111111111111" when X = 157 AND Y = 71 else
"111111111111" when X = 158 AND Y = 71 else
"111111111111" when X = 159 AND Y = 71 else
"111111111111" when X = 160 AND Y = 71 else
"111111111111" when X = 161 AND Y = 71 else
"111111111111" when X = 162 AND Y = 71 else
"111111111111" when X = 163 AND Y = 71 else
"111111111111" when X = 164 AND Y = 71 else
"111111111111" when X = 165 AND Y = 71 else
"111111111111" when X = 166 AND Y = 71 else
"111111111111" when X = 167 AND Y = 71 else
"111111111111" when X = 168 AND Y = 71 else
"111111111111" when X = 169 AND Y = 71 else
"111111111111" when X = 170 AND Y = 71 else
"111111111111" when X = 171 AND Y = 71 else
"111111111111" when X = 172 AND Y = 71 else
"111111111111" when X = 173 AND Y = 71 else
"111111111111" when X = 174 AND Y = 71 else
"111111111111" when X = 175 AND Y = 71 else
"111111111111" when X = 176 AND Y = 71 else
"111111111111" when X = 177 AND Y = 71 else
"111111111111" when X = 178 AND Y = 71 else
"111111111111" when X = 179 AND Y = 71 else
"111111111111" when X = 180 AND Y = 71 else
"111111111111" when X = 181 AND Y = 71 else
"111111111111" when X = 182 AND Y = 71 else
"111111111111" when X = 183 AND Y = 71 else
"111111111111" when X = 184 AND Y = 71 else
"111111111111" when X = 185 AND Y = 71 else
"111111111111" when X = 186 AND Y = 71 else
"111111111111" when X = 187 AND Y = 71 else
"111111111111" when X = 188 AND Y = 71 else
"111111111111" when X = 189 AND Y = 71 else
"111111111111" when X = 190 AND Y = 71 else
"111111111111" when X = 191 AND Y = 71 else
"111111111111" when X = 192 AND Y = 71 else
"111111111111" when X = 193 AND Y = 71 else
"111111111111" when X = 194 AND Y = 71 else
"111111111111" when X = 195 AND Y = 71 else
"111111111111" when X = 196 AND Y = 71 else
"111111111111" when X = 197 AND Y = 71 else
"111111111111" when X = 198 AND Y = 71 else
"111111111111" when X = 199 AND Y = 71 else
"111111111111" when X = 200 AND Y = 71 else
"111111111111" when X = 201 AND Y = 71 else
"111111111111" when X = 202 AND Y = 71 else
"111111111111" when X = 203 AND Y = 71 else
"111111111111" when X = 204 AND Y = 71 else
"111111111111" when X = 205 AND Y = 71 else
"111111111111" when X = 206 AND Y = 71 else
"111111111111" when X = 207 AND Y = 71 else
"111111111111" when X = 208 AND Y = 71 else
"111111111111" when X = 209 AND Y = 71 else
"111111111111" when X = 210 AND Y = 71 else
"111111111111" when X = 211 AND Y = 71 else
"111111111111" when X = 212 AND Y = 71 else
"111111111111" when X = 213 AND Y = 71 else
"111111111111" when X = 214 AND Y = 71 else
"111111111111" when X = 215 AND Y = 71 else
"111111111111" when X = 216 AND Y = 71 else
"111111111111" when X = 217 AND Y = 71 else
"111111111111" when X = 218 AND Y = 71 else
"111111111111" when X = 219 AND Y = 71 else
"111111111111" when X = 220 AND Y = 71 else
"111111111111" when X = 221 AND Y = 71 else
"111111111111" when X = 222 AND Y = 71 else
"111111111111" when X = 223 AND Y = 71 else
"111111111111" when X = 224 AND Y = 71 else
"111111111111" when X = 225 AND Y = 71 else
"111111111111" when X = 226 AND Y = 71 else
"111111111111" when X = 227 AND Y = 71 else
"111111111111" when X = 228 AND Y = 71 else
"111111111111" when X = 229 AND Y = 71 else
"111111111111" when X = 230 AND Y = 71 else
"111111111111" when X = 231 AND Y = 71 else
"111111111111" when X = 232 AND Y = 71 else
"111111111111" when X = 233 AND Y = 71 else
"111111111111" when X = 234 AND Y = 71 else
"111111111111" when X = 235 AND Y = 71 else
"111111111111" when X = 236 AND Y = 71 else
"111111111111" when X = 237 AND Y = 71 else
"111111111111" when X = 238 AND Y = 71 else
"111111111111" when X = 239 AND Y = 71 else
"111111111111" when X = 240 AND Y = 71 else
"111111111111" when X = 241 AND Y = 71 else
"111111111111" when X = 242 AND Y = 71 else
"111111111111" when X = 243 AND Y = 71 else
"111111111111" when X = 244 AND Y = 71 else
"111111111111" when X = 245 AND Y = 71 else
"111111111111" when X = 246 AND Y = 71 else
"111111111111" when X = 247 AND Y = 71 else
"111111111111" when X = 248 AND Y = 71 else
"111111111111" when X = 249 AND Y = 71 else
"111111111111" when X = 250 AND Y = 71 else
"111111111111" when X = 251 AND Y = 71 else
"111111111111" when X = 252 AND Y = 71 else
"111111111111" when X = 253 AND Y = 71 else
"111111111111" when X = 254 AND Y = 71 else
"111111111111" when X = 255 AND Y = 71 else
"111111111111" when X = 256 AND Y = 71 else
"111111111111" when X = 257 AND Y = 71 else
"111111111111" when X = 258 AND Y = 71 else
"111111111111" when X = 259 AND Y = 71 else
"111111111111" when X = 260 AND Y = 71 else
"111111111111" when X = 261 AND Y = 71 else
"111111111111" when X = 262 AND Y = 71 else
"111111111111" when X = 263 AND Y = 71 else
"111111111111" when X = 264 AND Y = 71 else
"110111011111" when X = 265 AND Y = 71 else
"110111011111" when X = 266 AND Y = 71 else
"110111011111" when X = 267 AND Y = 71 else
"110111011111" when X = 268 AND Y = 71 else
"110111011111" when X = 269 AND Y = 71 else
"110111011111" when X = 270 AND Y = 71 else
"110111011111" when X = 271 AND Y = 71 else
"110111011111" when X = 272 AND Y = 71 else
"110111011111" when X = 273 AND Y = 71 else
"110111011111" when X = 274 AND Y = 71 else
"110111011111" when X = 275 AND Y = 71 else
"110111011111" when X = 276 AND Y = 71 else
"110111011111" when X = 277 AND Y = 71 else
"110111011111" when X = 278 AND Y = 71 else
"110111011111" when X = 279 AND Y = 71 else
"000000000000" when X = 280 AND Y = 71 else
"000000000000" when X = 281 AND Y = 71 else
"000000000000" when X = 282 AND Y = 71 else
"000000000000" when X = 283 AND Y = 71 else
"000000000000" when X = 284 AND Y = 71 else
"000000000000" when X = 285 AND Y = 71 else
"000000000000" when X = 286 AND Y = 71 else
"000000000000" when X = 287 AND Y = 71 else
"000000000000" when X = 288 AND Y = 71 else
"000000000000" when X = 289 AND Y = 71 else
"000000000000" when X = 290 AND Y = 71 else
"000000000000" when X = 291 AND Y = 71 else
"000000000000" when X = 292 AND Y = 71 else
"000000000000" when X = 293 AND Y = 71 else
"000000000000" when X = 294 AND Y = 71 else
"000000000000" when X = 295 AND Y = 71 else
"000000000000" when X = 296 AND Y = 71 else
"000000000000" when X = 297 AND Y = 71 else
"000000000000" when X = 298 AND Y = 71 else
"000000000000" when X = 299 AND Y = 71 else
"000000000000" when X = 300 AND Y = 71 else
"000000000000" when X = 301 AND Y = 71 else
"000000000000" when X = 302 AND Y = 71 else
"000000000000" when X = 303 AND Y = 71 else
"000000000000" when X = 304 AND Y = 71 else
"000000000000" when X = 305 AND Y = 71 else
"000000000000" when X = 306 AND Y = 71 else
"000000000000" when X = 307 AND Y = 71 else
"000000000000" when X = 308 AND Y = 71 else
"000000000000" when X = 309 AND Y = 71 else
"000000000000" when X = 310 AND Y = 71 else
"000000000000" when X = 311 AND Y = 71 else
"000000000000" when X = 312 AND Y = 71 else
"000000000000" when X = 313 AND Y = 71 else
"000000000000" when X = 314 AND Y = 71 else
"000000000000" when X = 315 AND Y = 71 else
"000000000000" when X = 316 AND Y = 71 else
"000000000000" when X = 317 AND Y = 71 else
"000000000000" when X = 318 AND Y = 71 else
"000000000000" when X = 319 AND Y = 71 else
"000000000000" when X = 320 AND Y = 71 else
"000000000000" when X = 321 AND Y = 71 else
"000000000000" when X = 322 AND Y = 71 else
"000000000000" when X = 323 AND Y = 71 else
"000000000000" when X = 324 AND Y = 71 else
"100010011101" when X = 0 AND Y = 72 else
"100010011101" when X = 1 AND Y = 72 else
"100010011101" when X = 2 AND Y = 72 else
"100010011101" when X = 3 AND Y = 72 else
"100010011101" when X = 4 AND Y = 72 else
"100010011101" when X = 5 AND Y = 72 else
"100010011101" when X = 6 AND Y = 72 else
"100010011101" when X = 7 AND Y = 72 else
"100010011101" when X = 8 AND Y = 72 else
"100010011101" when X = 9 AND Y = 72 else
"100010011101" when X = 10 AND Y = 72 else
"100010011101" when X = 11 AND Y = 72 else
"100010011101" when X = 12 AND Y = 72 else
"100010011101" when X = 13 AND Y = 72 else
"100010011101" when X = 14 AND Y = 72 else
"100010011101" when X = 15 AND Y = 72 else
"100010011101" when X = 16 AND Y = 72 else
"100010011101" when X = 17 AND Y = 72 else
"100010011101" when X = 18 AND Y = 72 else
"100010011101" when X = 19 AND Y = 72 else
"100010011101" when X = 20 AND Y = 72 else
"100010011101" when X = 21 AND Y = 72 else
"100010011101" when X = 22 AND Y = 72 else
"100010011101" when X = 23 AND Y = 72 else
"100010011101" when X = 24 AND Y = 72 else
"100010011101" when X = 25 AND Y = 72 else
"100010011101" when X = 26 AND Y = 72 else
"100010011101" when X = 27 AND Y = 72 else
"100010011101" when X = 28 AND Y = 72 else
"100010011101" when X = 29 AND Y = 72 else
"110111011111" when X = 30 AND Y = 72 else
"110111011111" when X = 31 AND Y = 72 else
"110111011111" when X = 32 AND Y = 72 else
"110111011111" when X = 33 AND Y = 72 else
"110111011111" when X = 34 AND Y = 72 else
"110111011111" when X = 35 AND Y = 72 else
"110111011111" when X = 36 AND Y = 72 else
"110111011111" when X = 37 AND Y = 72 else
"110111011111" when X = 38 AND Y = 72 else
"110111011111" when X = 39 AND Y = 72 else
"110111011111" when X = 40 AND Y = 72 else
"110111011111" when X = 41 AND Y = 72 else
"110111011111" when X = 42 AND Y = 72 else
"110111011111" when X = 43 AND Y = 72 else
"110111011111" when X = 44 AND Y = 72 else
"110111011111" when X = 45 AND Y = 72 else
"110111011111" when X = 46 AND Y = 72 else
"110111011111" when X = 47 AND Y = 72 else
"110111011111" when X = 48 AND Y = 72 else
"110111011111" when X = 49 AND Y = 72 else
"110111011111" when X = 50 AND Y = 72 else
"110111011111" when X = 51 AND Y = 72 else
"110111011111" when X = 52 AND Y = 72 else
"110111011111" when X = 53 AND Y = 72 else
"110111011111" when X = 54 AND Y = 72 else
"110111011111" when X = 55 AND Y = 72 else
"110111011111" when X = 56 AND Y = 72 else
"110111011111" when X = 57 AND Y = 72 else
"110111011111" when X = 58 AND Y = 72 else
"110111011111" when X = 59 AND Y = 72 else
"110111011111" when X = 60 AND Y = 72 else
"110111011111" when X = 61 AND Y = 72 else
"110111011111" when X = 62 AND Y = 72 else
"110111011111" when X = 63 AND Y = 72 else
"110111011111" when X = 64 AND Y = 72 else
"110111011111" when X = 65 AND Y = 72 else
"110111011111" when X = 66 AND Y = 72 else
"110111011111" when X = 67 AND Y = 72 else
"110111011111" when X = 68 AND Y = 72 else
"110111011111" when X = 69 AND Y = 72 else
"110111011111" when X = 70 AND Y = 72 else
"110111011111" when X = 71 AND Y = 72 else
"110111011111" when X = 72 AND Y = 72 else
"110111011111" when X = 73 AND Y = 72 else
"110111011111" when X = 74 AND Y = 72 else
"110111011111" when X = 75 AND Y = 72 else
"110111011111" when X = 76 AND Y = 72 else
"110111011111" when X = 77 AND Y = 72 else
"110111011111" when X = 78 AND Y = 72 else
"110111011111" when X = 79 AND Y = 72 else
"110111011111" when X = 80 AND Y = 72 else
"110111011111" when X = 81 AND Y = 72 else
"110111011111" when X = 82 AND Y = 72 else
"110111011111" when X = 83 AND Y = 72 else
"110111011111" when X = 84 AND Y = 72 else
"110111011111" when X = 85 AND Y = 72 else
"110111011111" when X = 86 AND Y = 72 else
"110111011111" when X = 87 AND Y = 72 else
"110111011111" when X = 88 AND Y = 72 else
"110111011111" when X = 89 AND Y = 72 else
"110111011111" when X = 90 AND Y = 72 else
"110111011111" when X = 91 AND Y = 72 else
"110111011111" when X = 92 AND Y = 72 else
"110111011111" when X = 93 AND Y = 72 else
"110111011111" when X = 94 AND Y = 72 else
"110111011111" when X = 95 AND Y = 72 else
"110111011111" when X = 96 AND Y = 72 else
"110111011111" when X = 97 AND Y = 72 else
"110111011111" when X = 98 AND Y = 72 else
"110111011111" when X = 99 AND Y = 72 else
"110111011111" when X = 100 AND Y = 72 else
"110111011111" when X = 101 AND Y = 72 else
"110111011111" when X = 102 AND Y = 72 else
"110111011111" when X = 103 AND Y = 72 else
"110111011111" when X = 104 AND Y = 72 else
"111111111111" when X = 105 AND Y = 72 else
"111111111111" when X = 106 AND Y = 72 else
"111111111111" when X = 107 AND Y = 72 else
"111111111111" when X = 108 AND Y = 72 else
"111111111111" when X = 109 AND Y = 72 else
"111111111111" when X = 110 AND Y = 72 else
"111111111111" when X = 111 AND Y = 72 else
"111111111111" when X = 112 AND Y = 72 else
"111111111111" when X = 113 AND Y = 72 else
"111111111111" when X = 114 AND Y = 72 else
"111111111111" when X = 115 AND Y = 72 else
"111111111111" when X = 116 AND Y = 72 else
"111111111111" when X = 117 AND Y = 72 else
"111111111111" when X = 118 AND Y = 72 else
"111111111111" when X = 119 AND Y = 72 else
"111111111111" when X = 120 AND Y = 72 else
"111111111111" when X = 121 AND Y = 72 else
"111111111111" when X = 122 AND Y = 72 else
"111111111111" when X = 123 AND Y = 72 else
"111111111111" when X = 124 AND Y = 72 else
"111111111111" when X = 125 AND Y = 72 else
"111111111111" when X = 126 AND Y = 72 else
"111111111111" when X = 127 AND Y = 72 else
"111111111111" when X = 128 AND Y = 72 else
"111111111111" when X = 129 AND Y = 72 else
"111111111111" when X = 130 AND Y = 72 else
"111111111111" when X = 131 AND Y = 72 else
"111111111111" when X = 132 AND Y = 72 else
"111111111111" when X = 133 AND Y = 72 else
"111111111111" when X = 134 AND Y = 72 else
"111111111111" when X = 135 AND Y = 72 else
"111111111111" when X = 136 AND Y = 72 else
"111111111111" when X = 137 AND Y = 72 else
"111111111111" when X = 138 AND Y = 72 else
"111111111111" when X = 139 AND Y = 72 else
"111111111111" when X = 140 AND Y = 72 else
"111111111111" when X = 141 AND Y = 72 else
"111111111111" when X = 142 AND Y = 72 else
"111111111111" when X = 143 AND Y = 72 else
"111111111111" when X = 144 AND Y = 72 else
"111111111111" when X = 145 AND Y = 72 else
"111111111111" when X = 146 AND Y = 72 else
"111111111111" when X = 147 AND Y = 72 else
"111111111111" when X = 148 AND Y = 72 else
"111111111111" when X = 149 AND Y = 72 else
"111111111111" when X = 150 AND Y = 72 else
"111111111111" when X = 151 AND Y = 72 else
"111111111111" when X = 152 AND Y = 72 else
"111111111111" when X = 153 AND Y = 72 else
"111111111111" when X = 154 AND Y = 72 else
"111111111111" when X = 155 AND Y = 72 else
"111111111111" when X = 156 AND Y = 72 else
"111111111111" when X = 157 AND Y = 72 else
"111111111111" when X = 158 AND Y = 72 else
"111111111111" when X = 159 AND Y = 72 else
"111111111111" when X = 160 AND Y = 72 else
"111111111111" when X = 161 AND Y = 72 else
"111111111111" when X = 162 AND Y = 72 else
"111111111111" when X = 163 AND Y = 72 else
"111111111111" when X = 164 AND Y = 72 else
"111111111111" when X = 165 AND Y = 72 else
"111111111111" when X = 166 AND Y = 72 else
"111111111111" when X = 167 AND Y = 72 else
"111111111111" when X = 168 AND Y = 72 else
"111111111111" when X = 169 AND Y = 72 else
"111111111111" when X = 170 AND Y = 72 else
"111111111111" when X = 171 AND Y = 72 else
"111111111111" when X = 172 AND Y = 72 else
"111111111111" when X = 173 AND Y = 72 else
"111111111111" when X = 174 AND Y = 72 else
"111111111111" when X = 175 AND Y = 72 else
"111111111111" when X = 176 AND Y = 72 else
"111111111111" when X = 177 AND Y = 72 else
"111111111111" when X = 178 AND Y = 72 else
"111111111111" when X = 179 AND Y = 72 else
"111111111111" when X = 180 AND Y = 72 else
"111111111111" when X = 181 AND Y = 72 else
"111111111111" when X = 182 AND Y = 72 else
"111111111111" when X = 183 AND Y = 72 else
"111111111111" when X = 184 AND Y = 72 else
"111111111111" when X = 185 AND Y = 72 else
"111111111111" when X = 186 AND Y = 72 else
"111111111111" when X = 187 AND Y = 72 else
"111111111111" when X = 188 AND Y = 72 else
"111111111111" when X = 189 AND Y = 72 else
"111111111111" when X = 190 AND Y = 72 else
"111111111111" when X = 191 AND Y = 72 else
"111111111111" when X = 192 AND Y = 72 else
"111111111111" when X = 193 AND Y = 72 else
"111111111111" when X = 194 AND Y = 72 else
"111111111111" when X = 195 AND Y = 72 else
"111111111111" when X = 196 AND Y = 72 else
"111111111111" when X = 197 AND Y = 72 else
"111111111111" when X = 198 AND Y = 72 else
"111111111111" when X = 199 AND Y = 72 else
"111111111111" when X = 200 AND Y = 72 else
"111111111111" when X = 201 AND Y = 72 else
"111111111111" when X = 202 AND Y = 72 else
"111111111111" when X = 203 AND Y = 72 else
"111111111111" when X = 204 AND Y = 72 else
"111111111111" when X = 205 AND Y = 72 else
"111111111111" when X = 206 AND Y = 72 else
"111111111111" when X = 207 AND Y = 72 else
"111111111111" when X = 208 AND Y = 72 else
"111111111111" when X = 209 AND Y = 72 else
"111111111111" when X = 210 AND Y = 72 else
"111111111111" when X = 211 AND Y = 72 else
"111111111111" when X = 212 AND Y = 72 else
"111111111111" when X = 213 AND Y = 72 else
"111111111111" when X = 214 AND Y = 72 else
"111111111111" when X = 215 AND Y = 72 else
"111111111111" when X = 216 AND Y = 72 else
"111111111111" when X = 217 AND Y = 72 else
"111111111111" when X = 218 AND Y = 72 else
"111111111111" when X = 219 AND Y = 72 else
"111111111111" when X = 220 AND Y = 72 else
"111111111111" when X = 221 AND Y = 72 else
"111111111111" when X = 222 AND Y = 72 else
"111111111111" when X = 223 AND Y = 72 else
"111111111111" when X = 224 AND Y = 72 else
"111111111111" when X = 225 AND Y = 72 else
"111111111111" when X = 226 AND Y = 72 else
"111111111111" when X = 227 AND Y = 72 else
"111111111111" when X = 228 AND Y = 72 else
"111111111111" when X = 229 AND Y = 72 else
"111111111111" when X = 230 AND Y = 72 else
"111111111111" when X = 231 AND Y = 72 else
"111111111111" when X = 232 AND Y = 72 else
"111111111111" when X = 233 AND Y = 72 else
"111111111111" when X = 234 AND Y = 72 else
"111111111111" when X = 235 AND Y = 72 else
"111111111111" when X = 236 AND Y = 72 else
"111111111111" when X = 237 AND Y = 72 else
"111111111111" when X = 238 AND Y = 72 else
"111111111111" when X = 239 AND Y = 72 else
"111111111111" when X = 240 AND Y = 72 else
"111111111111" when X = 241 AND Y = 72 else
"111111111111" when X = 242 AND Y = 72 else
"111111111111" when X = 243 AND Y = 72 else
"111111111111" when X = 244 AND Y = 72 else
"111111111111" when X = 245 AND Y = 72 else
"111111111111" when X = 246 AND Y = 72 else
"111111111111" when X = 247 AND Y = 72 else
"111111111111" when X = 248 AND Y = 72 else
"111111111111" when X = 249 AND Y = 72 else
"111111111111" when X = 250 AND Y = 72 else
"111111111111" when X = 251 AND Y = 72 else
"111111111111" when X = 252 AND Y = 72 else
"111111111111" when X = 253 AND Y = 72 else
"111111111111" when X = 254 AND Y = 72 else
"111111111111" when X = 255 AND Y = 72 else
"111111111111" when X = 256 AND Y = 72 else
"111111111111" when X = 257 AND Y = 72 else
"111111111111" when X = 258 AND Y = 72 else
"111111111111" when X = 259 AND Y = 72 else
"111111111111" when X = 260 AND Y = 72 else
"111111111111" when X = 261 AND Y = 72 else
"111111111111" when X = 262 AND Y = 72 else
"111111111111" when X = 263 AND Y = 72 else
"111111111111" when X = 264 AND Y = 72 else
"110111011111" when X = 265 AND Y = 72 else
"110111011111" when X = 266 AND Y = 72 else
"110111011111" when X = 267 AND Y = 72 else
"110111011111" when X = 268 AND Y = 72 else
"110111011111" when X = 269 AND Y = 72 else
"110111011111" when X = 270 AND Y = 72 else
"110111011111" when X = 271 AND Y = 72 else
"110111011111" when X = 272 AND Y = 72 else
"110111011111" when X = 273 AND Y = 72 else
"110111011111" when X = 274 AND Y = 72 else
"110111011111" when X = 275 AND Y = 72 else
"110111011111" when X = 276 AND Y = 72 else
"110111011111" when X = 277 AND Y = 72 else
"110111011111" when X = 278 AND Y = 72 else
"110111011111" when X = 279 AND Y = 72 else
"000000000000" when X = 280 AND Y = 72 else
"000000000000" when X = 281 AND Y = 72 else
"000000000000" when X = 282 AND Y = 72 else
"000000000000" when X = 283 AND Y = 72 else
"000000000000" when X = 284 AND Y = 72 else
"000000000000" when X = 285 AND Y = 72 else
"000000000000" when X = 286 AND Y = 72 else
"000000000000" when X = 287 AND Y = 72 else
"000000000000" when X = 288 AND Y = 72 else
"000000000000" when X = 289 AND Y = 72 else
"000000000000" when X = 290 AND Y = 72 else
"000000000000" when X = 291 AND Y = 72 else
"000000000000" when X = 292 AND Y = 72 else
"000000000000" when X = 293 AND Y = 72 else
"000000000000" when X = 294 AND Y = 72 else
"000000000000" when X = 295 AND Y = 72 else
"000000000000" when X = 296 AND Y = 72 else
"000000000000" when X = 297 AND Y = 72 else
"000000000000" when X = 298 AND Y = 72 else
"000000000000" when X = 299 AND Y = 72 else
"000000000000" when X = 300 AND Y = 72 else
"000000000000" when X = 301 AND Y = 72 else
"000000000000" when X = 302 AND Y = 72 else
"000000000000" when X = 303 AND Y = 72 else
"000000000000" when X = 304 AND Y = 72 else
"000000000000" when X = 305 AND Y = 72 else
"000000000000" when X = 306 AND Y = 72 else
"000000000000" when X = 307 AND Y = 72 else
"000000000000" when X = 308 AND Y = 72 else
"000000000000" when X = 309 AND Y = 72 else
"000000000000" when X = 310 AND Y = 72 else
"000000000000" when X = 311 AND Y = 72 else
"000000000000" when X = 312 AND Y = 72 else
"000000000000" when X = 313 AND Y = 72 else
"000000000000" when X = 314 AND Y = 72 else
"000000000000" when X = 315 AND Y = 72 else
"000000000000" when X = 316 AND Y = 72 else
"000000000000" when X = 317 AND Y = 72 else
"000000000000" when X = 318 AND Y = 72 else
"000000000000" when X = 319 AND Y = 72 else
"000000000000" when X = 320 AND Y = 72 else
"000000000000" when X = 321 AND Y = 72 else
"000000000000" when X = 322 AND Y = 72 else
"000000000000" when X = 323 AND Y = 72 else
"000000000000" when X = 324 AND Y = 72 else
"100010011101" when X = 0 AND Y = 73 else
"100010011101" when X = 1 AND Y = 73 else
"100010011101" when X = 2 AND Y = 73 else
"100010011101" when X = 3 AND Y = 73 else
"100010011101" when X = 4 AND Y = 73 else
"100010011101" when X = 5 AND Y = 73 else
"100010011101" when X = 6 AND Y = 73 else
"100010011101" when X = 7 AND Y = 73 else
"100010011101" when X = 8 AND Y = 73 else
"100010011101" when X = 9 AND Y = 73 else
"100010011101" when X = 10 AND Y = 73 else
"100010011101" when X = 11 AND Y = 73 else
"100010011101" when X = 12 AND Y = 73 else
"100010011101" when X = 13 AND Y = 73 else
"100010011101" when X = 14 AND Y = 73 else
"100010011101" when X = 15 AND Y = 73 else
"100010011101" when X = 16 AND Y = 73 else
"100010011101" when X = 17 AND Y = 73 else
"100010011101" when X = 18 AND Y = 73 else
"100010011101" when X = 19 AND Y = 73 else
"100010011101" when X = 20 AND Y = 73 else
"100010011101" when X = 21 AND Y = 73 else
"100010011101" when X = 22 AND Y = 73 else
"100010011101" when X = 23 AND Y = 73 else
"100010011101" when X = 24 AND Y = 73 else
"100010011101" when X = 25 AND Y = 73 else
"100010011101" when X = 26 AND Y = 73 else
"100010011101" when X = 27 AND Y = 73 else
"100010011101" when X = 28 AND Y = 73 else
"100010011101" when X = 29 AND Y = 73 else
"110111011111" when X = 30 AND Y = 73 else
"110111011111" when X = 31 AND Y = 73 else
"110111011111" when X = 32 AND Y = 73 else
"110111011111" when X = 33 AND Y = 73 else
"110111011111" when X = 34 AND Y = 73 else
"110111011111" when X = 35 AND Y = 73 else
"110111011111" when X = 36 AND Y = 73 else
"110111011111" when X = 37 AND Y = 73 else
"110111011111" when X = 38 AND Y = 73 else
"110111011111" when X = 39 AND Y = 73 else
"110111011111" when X = 40 AND Y = 73 else
"110111011111" when X = 41 AND Y = 73 else
"110111011111" when X = 42 AND Y = 73 else
"110111011111" when X = 43 AND Y = 73 else
"110111011111" when X = 44 AND Y = 73 else
"110111011111" when X = 45 AND Y = 73 else
"110111011111" when X = 46 AND Y = 73 else
"110111011111" when X = 47 AND Y = 73 else
"110111011111" when X = 48 AND Y = 73 else
"110111011111" when X = 49 AND Y = 73 else
"110111011111" when X = 50 AND Y = 73 else
"110111011111" when X = 51 AND Y = 73 else
"110111011111" when X = 52 AND Y = 73 else
"110111011111" when X = 53 AND Y = 73 else
"110111011111" when X = 54 AND Y = 73 else
"110111011111" when X = 55 AND Y = 73 else
"110111011111" when X = 56 AND Y = 73 else
"110111011111" when X = 57 AND Y = 73 else
"110111011111" when X = 58 AND Y = 73 else
"110111011111" when X = 59 AND Y = 73 else
"110111011111" when X = 60 AND Y = 73 else
"110111011111" when X = 61 AND Y = 73 else
"110111011111" when X = 62 AND Y = 73 else
"110111011111" when X = 63 AND Y = 73 else
"110111011111" when X = 64 AND Y = 73 else
"110111011111" when X = 65 AND Y = 73 else
"110111011111" when X = 66 AND Y = 73 else
"110111011111" when X = 67 AND Y = 73 else
"110111011111" when X = 68 AND Y = 73 else
"110111011111" when X = 69 AND Y = 73 else
"110111011111" when X = 70 AND Y = 73 else
"110111011111" when X = 71 AND Y = 73 else
"110111011111" when X = 72 AND Y = 73 else
"110111011111" when X = 73 AND Y = 73 else
"110111011111" when X = 74 AND Y = 73 else
"110111011111" when X = 75 AND Y = 73 else
"110111011111" when X = 76 AND Y = 73 else
"110111011111" when X = 77 AND Y = 73 else
"110111011111" when X = 78 AND Y = 73 else
"110111011111" when X = 79 AND Y = 73 else
"110111011111" when X = 80 AND Y = 73 else
"110111011111" when X = 81 AND Y = 73 else
"110111011111" when X = 82 AND Y = 73 else
"110111011111" when X = 83 AND Y = 73 else
"110111011111" when X = 84 AND Y = 73 else
"110111011111" when X = 85 AND Y = 73 else
"110111011111" when X = 86 AND Y = 73 else
"110111011111" when X = 87 AND Y = 73 else
"110111011111" when X = 88 AND Y = 73 else
"110111011111" when X = 89 AND Y = 73 else
"110111011111" when X = 90 AND Y = 73 else
"110111011111" when X = 91 AND Y = 73 else
"110111011111" when X = 92 AND Y = 73 else
"110111011111" when X = 93 AND Y = 73 else
"110111011111" when X = 94 AND Y = 73 else
"110111011111" when X = 95 AND Y = 73 else
"110111011111" when X = 96 AND Y = 73 else
"110111011111" when X = 97 AND Y = 73 else
"110111011111" when X = 98 AND Y = 73 else
"110111011111" when X = 99 AND Y = 73 else
"110111011111" when X = 100 AND Y = 73 else
"110111011111" when X = 101 AND Y = 73 else
"110111011111" when X = 102 AND Y = 73 else
"110111011111" when X = 103 AND Y = 73 else
"110111011111" when X = 104 AND Y = 73 else
"111111111111" when X = 105 AND Y = 73 else
"111111111111" when X = 106 AND Y = 73 else
"111111111111" when X = 107 AND Y = 73 else
"111111111111" when X = 108 AND Y = 73 else
"111111111111" when X = 109 AND Y = 73 else
"111111111111" when X = 110 AND Y = 73 else
"111111111111" when X = 111 AND Y = 73 else
"111111111111" when X = 112 AND Y = 73 else
"111111111111" when X = 113 AND Y = 73 else
"111111111111" when X = 114 AND Y = 73 else
"111111111111" when X = 115 AND Y = 73 else
"111111111111" when X = 116 AND Y = 73 else
"111111111111" when X = 117 AND Y = 73 else
"111111111111" when X = 118 AND Y = 73 else
"111111111111" when X = 119 AND Y = 73 else
"111111111111" when X = 120 AND Y = 73 else
"111111111111" when X = 121 AND Y = 73 else
"111111111111" when X = 122 AND Y = 73 else
"111111111111" when X = 123 AND Y = 73 else
"111111111111" when X = 124 AND Y = 73 else
"111111111111" when X = 125 AND Y = 73 else
"111111111111" when X = 126 AND Y = 73 else
"111111111111" when X = 127 AND Y = 73 else
"111111111111" when X = 128 AND Y = 73 else
"111111111111" when X = 129 AND Y = 73 else
"111111111111" when X = 130 AND Y = 73 else
"111111111111" when X = 131 AND Y = 73 else
"111111111111" when X = 132 AND Y = 73 else
"111111111111" when X = 133 AND Y = 73 else
"111111111111" when X = 134 AND Y = 73 else
"111111111111" when X = 135 AND Y = 73 else
"111111111111" when X = 136 AND Y = 73 else
"111111111111" when X = 137 AND Y = 73 else
"111111111111" when X = 138 AND Y = 73 else
"111111111111" when X = 139 AND Y = 73 else
"111111111111" when X = 140 AND Y = 73 else
"111111111111" when X = 141 AND Y = 73 else
"111111111111" when X = 142 AND Y = 73 else
"111111111111" when X = 143 AND Y = 73 else
"111111111111" when X = 144 AND Y = 73 else
"111111111111" when X = 145 AND Y = 73 else
"111111111111" when X = 146 AND Y = 73 else
"111111111111" when X = 147 AND Y = 73 else
"111111111111" when X = 148 AND Y = 73 else
"111111111111" when X = 149 AND Y = 73 else
"111111111111" when X = 150 AND Y = 73 else
"111111111111" when X = 151 AND Y = 73 else
"111111111111" when X = 152 AND Y = 73 else
"111111111111" when X = 153 AND Y = 73 else
"111111111111" when X = 154 AND Y = 73 else
"111111111111" when X = 155 AND Y = 73 else
"111111111111" when X = 156 AND Y = 73 else
"111111111111" when X = 157 AND Y = 73 else
"111111111111" when X = 158 AND Y = 73 else
"111111111111" when X = 159 AND Y = 73 else
"111111111111" when X = 160 AND Y = 73 else
"111111111111" when X = 161 AND Y = 73 else
"111111111111" when X = 162 AND Y = 73 else
"111111111111" when X = 163 AND Y = 73 else
"111111111111" when X = 164 AND Y = 73 else
"111111111111" when X = 165 AND Y = 73 else
"111111111111" when X = 166 AND Y = 73 else
"111111111111" when X = 167 AND Y = 73 else
"111111111111" when X = 168 AND Y = 73 else
"111111111111" when X = 169 AND Y = 73 else
"111111111111" when X = 170 AND Y = 73 else
"111111111111" when X = 171 AND Y = 73 else
"111111111111" when X = 172 AND Y = 73 else
"111111111111" when X = 173 AND Y = 73 else
"111111111111" when X = 174 AND Y = 73 else
"111111111111" when X = 175 AND Y = 73 else
"111111111111" when X = 176 AND Y = 73 else
"111111111111" when X = 177 AND Y = 73 else
"111111111111" when X = 178 AND Y = 73 else
"111111111111" when X = 179 AND Y = 73 else
"111111111111" when X = 180 AND Y = 73 else
"111111111111" when X = 181 AND Y = 73 else
"111111111111" when X = 182 AND Y = 73 else
"111111111111" when X = 183 AND Y = 73 else
"111111111111" when X = 184 AND Y = 73 else
"111111111111" when X = 185 AND Y = 73 else
"111111111111" when X = 186 AND Y = 73 else
"111111111111" when X = 187 AND Y = 73 else
"111111111111" when X = 188 AND Y = 73 else
"111111111111" when X = 189 AND Y = 73 else
"111111111111" when X = 190 AND Y = 73 else
"111111111111" when X = 191 AND Y = 73 else
"111111111111" when X = 192 AND Y = 73 else
"111111111111" when X = 193 AND Y = 73 else
"111111111111" when X = 194 AND Y = 73 else
"111111111111" when X = 195 AND Y = 73 else
"111111111111" when X = 196 AND Y = 73 else
"111111111111" when X = 197 AND Y = 73 else
"111111111111" when X = 198 AND Y = 73 else
"111111111111" when X = 199 AND Y = 73 else
"111111111111" when X = 200 AND Y = 73 else
"111111111111" when X = 201 AND Y = 73 else
"111111111111" when X = 202 AND Y = 73 else
"111111111111" when X = 203 AND Y = 73 else
"111111111111" when X = 204 AND Y = 73 else
"111111111111" when X = 205 AND Y = 73 else
"111111111111" when X = 206 AND Y = 73 else
"111111111111" when X = 207 AND Y = 73 else
"111111111111" when X = 208 AND Y = 73 else
"111111111111" when X = 209 AND Y = 73 else
"111111111111" when X = 210 AND Y = 73 else
"111111111111" when X = 211 AND Y = 73 else
"111111111111" when X = 212 AND Y = 73 else
"111111111111" when X = 213 AND Y = 73 else
"111111111111" when X = 214 AND Y = 73 else
"111111111111" when X = 215 AND Y = 73 else
"111111111111" when X = 216 AND Y = 73 else
"111111111111" when X = 217 AND Y = 73 else
"111111111111" when X = 218 AND Y = 73 else
"111111111111" when X = 219 AND Y = 73 else
"111111111111" when X = 220 AND Y = 73 else
"111111111111" when X = 221 AND Y = 73 else
"111111111111" when X = 222 AND Y = 73 else
"111111111111" when X = 223 AND Y = 73 else
"111111111111" when X = 224 AND Y = 73 else
"111111111111" when X = 225 AND Y = 73 else
"111111111111" when X = 226 AND Y = 73 else
"111111111111" when X = 227 AND Y = 73 else
"111111111111" when X = 228 AND Y = 73 else
"111111111111" when X = 229 AND Y = 73 else
"111111111111" when X = 230 AND Y = 73 else
"111111111111" when X = 231 AND Y = 73 else
"111111111111" when X = 232 AND Y = 73 else
"111111111111" when X = 233 AND Y = 73 else
"111111111111" when X = 234 AND Y = 73 else
"111111111111" when X = 235 AND Y = 73 else
"111111111111" when X = 236 AND Y = 73 else
"111111111111" when X = 237 AND Y = 73 else
"111111111111" when X = 238 AND Y = 73 else
"111111111111" when X = 239 AND Y = 73 else
"111111111111" when X = 240 AND Y = 73 else
"111111111111" when X = 241 AND Y = 73 else
"111111111111" when X = 242 AND Y = 73 else
"111111111111" when X = 243 AND Y = 73 else
"111111111111" when X = 244 AND Y = 73 else
"111111111111" when X = 245 AND Y = 73 else
"111111111111" when X = 246 AND Y = 73 else
"111111111111" when X = 247 AND Y = 73 else
"111111111111" when X = 248 AND Y = 73 else
"111111111111" when X = 249 AND Y = 73 else
"111111111111" when X = 250 AND Y = 73 else
"111111111111" when X = 251 AND Y = 73 else
"111111111111" when X = 252 AND Y = 73 else
"111111111111" when X = 253 AND Y = 73 else
"111111111111" when X = 254 AND Y = 73 else
"111111111111" when X = 255 AND Y = 73 else
"111111111111" when X = 256 AND Y = 73 else
"111111111111" when X = 257 AND Y = 73 else
"111111111111" when X = 258 AND Y = 73 else
"111111111111" when X = 259 AND Y = 73 else
"111111111111" when X = 260 AND Y = 73 else
"111111111111" when X = 261 AND Y = 73 else
"111111111111" when X = 262 AND Y = 73 else
"111111111111" when X = 263 AND Y = 73 else
"111111111111" when X = 264 AND Y = 73 else
"110111011111" when X = 265 AND Y = 73 else
"110111011111" when X = 266 AND Y = 73 else
"110111011111" when X = 267 AND Y = 73 else
"110111011111" when X = 268 AND Y = 73 else
"110111011111" when X = 269 AND Y = 73 else
"110111011111" when X = 270 AND Y = 73 else
"110111011111" when X = 271 AND Y = 73 else
"110111011111" when X = 272 AND Y = 73 else
"110111011111" when X = 273 AND Y = 73 else
"110111011111" when X = 274 AND Y = 73 else
"110111011111" when X = 275 AND Y = 73 else
"110111011111" when X = 276 AND Y = 73 else
"110111011111" when X = 277 AND Y = 73 else
"110111011111" when X = 278 AND Y = 73 else
"110111011111" when X = 279 AND Y = 73 else
"000000000000" when X = 280 AND Y = 73 else
"000000000000" when X = 281 AND Y = 73 else
"000000000000" when X = 282 AND Y = 73 else
"000000000000" when X = 283 AND Y = 73 else
"000000000000" when X = 284 AND Y = 73 else
"000000000000" when X = 285 AND Y = 73 else
"000000000000" when X = 286 AND Y = 73 else
"000000000000" when X = 287 AND Y = 73 else
"000000000000" when X = 288 AND Y = 73 else
"000000000000" when X = 289 AND Y = 73 else
"000000000000" when X = 290 AND Y = 73 else
"000000000000" when X = 291 AND Y = 73 else
"000000000000" when X = 292 AND Y = 73 else
"000000000000" when X = 293 AND Y = 73 else
"000000000000" when X = 294 AND Y = 73 else
"000000000000" when X = 295 AND Y = 73 else
"000000000000" when X = 296 AND Y = 73 else
"000000000000" when X = 297 AND Y = 73 else
"000000000000" when X = 298 AND Y = 73 else
"000000000000" when X = 299 AND Y = 73 else
"000000000000" when X = 300 AND Y = 73 else
"000000000000" when X = 301 AND Y = 73 else
"000000000000" when X = 302 AND Y = 73 else
"000000000000" when X = 303 AND Y = 73 else
"000000000000" when X = 304 AND Y = 73 else
"000000000000" when X = 305 AND Y = 73 else
"000000000000" when X = 306 AND Y = 73 else
"000000000000" when X = 307 AND Y = 73 else
"000000000000" when X = 308 AND Y = 73 else
"000000000000" when X = 309 AND Y = 73 else
"000000000000" when X = 310 AND Y = 73 else
"000000000000" when X = 311 AND Y = 73 else
"000000000000" when X = 312 AND Y = 73 else
"000000000000" when X = 313 AND Y = 73 else
"000000000000" when X = 314 AND Y = 73 else
"000000000000" when X = 315 AND Y = 73 else
"000000000000" when X = 316 AND Y = 73 else
"000000000000" when X = 317 AND Y = 73 else
"000000000000" when X = 318 AND Y = 73 else
"000000000000" when X = 319 AND Y = 73 else
"000000000000" when X = 320 AND Y = 73 else
"000000000000" when X = 321 AND Y = 73 else
"000000000000" when X = 322 AND Y = 73 else
"000000000000" when X = 323 AND Y = 73 else
"000000000000" when X = 324 AND Y = 73 else
"100010011101" when X = 0 AND Y = 74 else
"100010011101" when X = 1 AND Y = 74 else
"100010011101" when X = 2 AND Y = 74 else
"100010011101" when X = 3 AND Y = 74 else
"100010011101" when X = 4 AND Y = 74 else
"100010011101" when X = 5 AND Y = 74 else
"100010011101" when X = 6 AND Y = 74 else
"100010011101" when X = 7 AND Y = 74 else
"100010011101" when X = 8 AND Y = 74 else
"100010011101" when X = 9 AND Y = 74 else
"100010011101" when X = 10 AND Y = 74 else
"100010011101" when X = 11 AND Y = 74 else
"100010011101" when X = 12 AND Y = 74 else
"100010011101" when X = 13 AND Y = 74 else
"100010011101" when X = 14 AND Y = 74 else
"100010011101" when X = 15 AND Y = 74 else
"100010011101" when X = 16 AND Y = 74 else
"100010011101" when X = 17 AND Y = 74 else
"100010011101" when X = 18 AND Y = 74 else
"100010011101" when X = 19 AND Y = 74 else
"100010011101" when X = 20 AND Y = 74 else
"100010011101" when X = 21 AND Y = 74 else
"100010011101" when X = 22 AND Y = 74 else
"100010011101" when X = 23 AND Y = 74 else
"100010011101" when X = 24 AND Y = 74 else
"100010011101" when X = 25 AND Y = 74 else
"100010011101" when X = 26 AND Y = 74 else
"100010011101" when X = 27 AND Y = 74 else
"100010011101" when X = 28 AND Y = 74 else
"100010011101" when X = 29 AND Y = 74 else
"110111011111" when X = 30 AND Y = 74 else
"110111011111" when X = 31 AND Y = 74 else
"110111011111" when X = 32 AND Y = 74 else
"110111011111" when X = 33 AND Y = 74 else
"110111011111" when X = 34 AND Y = 74 else
"110111011111" when X = 35 AND Y = 74 else
"110111011111" when X = 36 AND Y = 74 else
"110111011111" when X = 37 AND Y = 74 else
"110111011111" when X = 38 AND Y = 74 else
"110111011111" when X = 39 AND Y = 74 else
"110111011111" when X = 40 AND Y = 74 else
"110111011111" when X = 41 AND Y = 74 else
"110111011111" when X = 42 AND Y = 74 else
"110111011111" when X = 43 AND Y = 74 else
"110111011111" when X = 44 AND Y = 74 else
"110111011111" when X = 45 AND Y = 74 else
"110111011111" when X = 46 AND Y = 74 else
"110111011111" when X = 47 AND Y = 74 else
"110111011111" when X = 48 AND Y = 74 else
"110111011111" when X = 49 AND Y = 74 else
"110111011111" when X = 50 AND Y = 74 else
"110111011111" when X = 51 AND Y = 74 else
"110111011111" when X = 52 AND Y = 74 else
"110111011111" when X = 53 AND Y = 74 else
"110111011111" when X = 54 AND Y = 74 else
"110111011111" when X = 55 AND Y = 74 else
"110111011111" when X = 56 AND Y = 74 else
"110111011111" when X = 57 AND Y = 74 else
"110111011111" when X = 58 AND Y = 74 else
"110111011111" when X = 59 AND Y = 74 else
"110111011111" when X = 60 AND Y = 74 else
"110111011111" when X = 61 AND Y = 74 else
"110111011111" when X = 62 AND Y = 74 else
"110111011111" when X = 63 AND Y = 74 else
"110111011111" when X = 64 AND Y = 74 else
"110111011111" when X = 65 AND Y = 74 else
"110111011111" when X = 66 AND Y = 74 else
"110111011111" when X = 67 AND Y = 74 else
"110111011111" when X = 68 AND Y = 74 else
"110111011111" when X = 69 AND Y = 74 else
"110111011111" when X = 70 AND Y = 74 else
"110111011111" when X = 71 AND Y = 74 else
"110111011111" when X = 72 AND Y = 74 else
"110111011111" when X = 73 AND Y = 74 else
"110111011111" when X = 74 AND Y = 74 else
"110111011111" when X = 75 AND Y = 74 else
"110111011111" when X = 76 AND Y = 74 else
"110111011111" when X = 77 AND Y = 74 else
"110111011111" when X = 78 AND Y = 74 else
"110111011111" when X = 79 AND Y = 74 else
"110111011111" when X = 80 AND Y = 74 else
"110111011111" when X = 81 AND Y = 74 else
"110111011111" when X = 82 AND Y = 74 else
"110111011111" when X = 83 AND Y = 74 else
"110111011111" when X = 84 AND Y = 74 else
"110111011111" when X = 85 AND Y = 74 else
"110111011111" when X = 86 AND Y = 74 else
"110111011111" when X = 87 AND Y = 74 else
"110111011111" when X = 88 AND Y = 74 else
"110111011111" when X = 89 AND Y = 74 else
"110111011111" when X = 90 AND Y = 74 else
"110111011111" when X = 91 AND Y = 74 else
"110111011111" when X = 92 AND Y = 74 else
"110111011111" when X = 93 AND Y = 74 else
"110111011111" when X = 94 AND Y = 74 else
"110111011111" when X = 95 AND Y = 74 else
"110111011111" when X = 96 AND Y = 74 else
"110111011111" when X = 97 AND Y = 74 else
"110111011111" when X = 98 AND Y = 74 else
"110111011111" when X = 99 AND Y = 74 else
"110111011111" when X = 100 AND Y = 74 else
"110111011111" when X = 101 AND Y = 74 else
"110111011111" when X = 102 AND Y = 74 else
"110111011111" when X = 103 AND Y = 74 else
"110111011111" when X = 104 AND Y = 74 else
"111111111111" when X = 105 AND Y = 74 else
"111111111111" when X = 106 AND Y = 74 else
"111111111111" when X = 107 AND Y = 74 else
"111111111111" when X = 108 AND Y = 74 else
"111111111111" when X = 109 AND Y = 74 else
"111111111111" when X = 110 AND Y = 74 else
"111111111111" when X = 111 AND Y = 74 else
"111111111111" when X = 112 AND Y = 74 else
"111111111111" when X = 113 AND Y = 74 else
"111111111111" when X = 114 AND Y = 74 else
"111111111111" when X = 115 AND Y = 74 else
"111111111111" when X = 116 AND Y = 74 else
"111111111111" when X = 117 AND Y = 74 else
"111111111111" when X = 118 AND Y = 74 else
"111111111111" when X = 119 AND Y = 74 else
"111111111111" when X = 120 AND Y = 74 else
"111111111111" when X = 121 AND Y = 74 else
"111111111111" when X = 122 AND Y = 74 else
"111111111111" when X = 123 AND Y = 74 else
"111111111111" when X = 124 AND Y = 74 else
"111111111111" when X = 125 AND Y = 74 else
"111111111111" when X = 126 AND Y = 74 else
"111111111111" when X = 127 AND Y = 74 else
"111111111111" when X = 128 AND Y = 74 else
"111111111111" when X = 129 AND Y = 74 else
"111111111111" when X = 130 AND Y = 74 else
"111111111111" when X = 131 AND Y = 74 else
"111111111111" when X = 132 AND Y = 74 else
"111111111111" when X = 133 AND Y = 74 else
"111111111111" when X = 134 AND Y = 74 else
"111111111111" when X = 135 AND Y = 74 else
"111111111111" when X = 136 AND Y = 74 else
"111111111111" when X = 137 AND Y = 74 else
"111111111111" when X = 138 AND Y = 74 else
"111111111111" when X = 139 AND Y = 74 else
"111111111111" when X = 140 AND Y = 74 else
"111111111111" when X = 141 AND Y = 74 else
"111111111111" when X = 142 AND Y = 74 else
"111111111111" when X = 143 AND Y = 74 else
"111111111111" when X = 144 AND Y = 74 else
"111111111111" when X = 145 AND Y = 74 else
"111111111111" when X = 146 AND Y = 74 else
"111111111111" when X = 147 AND Y = 74 else
"111111111111" when X = 148 AND Y = 74 else
"111111111111" when X = 149 AND Y = 74 else
"111111111111" when X = 150 AND Y = 74 else
"111111111111" when X = 151 AND Y = 74 else
"111111111111" when X = 152 AND Y = 74 else
"111111111111" when X = 153 AND Y = 74 else
"111111111111" when X = 154 AND Y = 74 else
"111111111111" when X = 155 AND Y = 74 else
"111111111111" when X = 156 AND Y = 74 else
"111111111111" when X = 157 AND Y = 74 else
"111111111111" when X = 158 AND Y = 74 else
"111111111111" when X = 159 AND Y = 74 else
"111111111111" when X = 160 AND Y = 74 else
"111111111111" when X = 161 AND Y = 74 else
"111111111111" when X = 162 AND Y = 74 else
"111111111111" when X = 163 AND Y = 74 else
"111111111111" when X = 164 AND Y = 74 else
"111111111111" when X = 165 AND Y = 74 else
"111111111111" when X = 166 AND Y = 74 else
"111111111111" when X = 167 AND Y = 74 else
"111111111111" when X = 168 AND Y = 74 else
"111111111111" when X = 169 AND Y = 74 else
"111111111111" when X = 170 AND Y = 74 else
"111111111111" when X = 171 AND Y = 74 else
"111111111111" when X = 172 AND Y = 74 else
"111111111111" when X = 173 AND Y = 74 else
"111111111111" when X = 174 AND Y = 74 else
"111111111111" when X = 175 AND Y = 74 else
"111111111111" when X = 176 AND Y = 74 else
"111111111111" when X = 177 AND Y = 74 else
"111111111111" when X = 178 AND Y = 74 else
"111111111111" when X = 179 AND Y = 74 else
"111111111111" when X = 180 AND Y = 74 else
"111111111111" when X = 181 AND Y = 74 else
"111111111111" when X = 182 AND Y = 74 else
"111111111111" when X = 183 AND Y = 74 else
"111111111111" when X = 184 AND Y = 74 else
"111111111111" when X = 185 AND Y = 74 else
"111111111111" when X = 186 AND Y = 74 else
"111111111111" when X = 187 AND Y = 74 else
"111111111111" when X = 188 AND Y = 74 else
"111111111111" when X = 189 AND Y = 74 else
"111111111111" when X = 190 AND Y = 74 else
"111111111111" when X = 191 AND Y = 74 else
"111111111111" when X = 192 AND Y = 74 else
"111111111111" when X = 193 AND Y = 74 else
"111111111111" when X = 194 AND Y = 74 else
"111111111111" when X = 195 AND Y = 74 else
"111111111111" when X = 196 AND Y = 74 else
"111111111111" when X = 197 AND Y = 74 else
"111111111111" when X = 198 AND Y = 74 else
"111111111111" when X = 199 AND Y = 74 else
"111111111111" when X = 200 AND Y = 74 else
"111111111111" when X = 201 AND Y = 74 else
"111111111111" when X = 202 AND Y = 74 else
"111111111111" when X = 203 AND Y = 74 else
"111111111111" when X = 204 AND Y = 74 else
"111111111111" when X = 205 AND Y = 74 else
"111111111111" when X = 206 AND Y = 74 else
"111111111111" when X = 207 AND Y = 74 else
"111111111111" when X = 208 AND Y = 74 else
"111111111111" when X = 209 AND Y = 74 else
"111111111111" when X = 210 AND Y = 74 else
"111111111111" when X = 211 AND Y = 74 else
"111111111111" when X = 212 AND Y = 74 else
"111111111111" when X = 213 AND Y = 74 else
"111111111111" when X = 214 AND Y = 74 else
"111111111111" when X = 215 AND Y = 74 else
"111111111111" when X = 216 AND Y = 74 else
"111111111111" when X = 217 AND Y = 74 else
"111111111111" when X = 218 AND Y = 74 else
"111111111111" when X = 219 AND Y = 74 else
"111111111111" when X = 220 AND Y = 74 else
"111111111111" when X = 221 AND Y = 74 else
"111111111111" when X = 222 AND Y = 74 else
"111111111111" when X = 223 AND Y = 74 else
"111111111111" when X = 224 AND Y = 74 else
"111111111111" when X = 225 AND Y = 74 else
"111111111111" when X = 226 AND Y = 74 else
"111111111111" when X = 227 AND Y = 74 else
"111111111111" when X = 228 AND Y = 74 else
"111111111111" when X = 229 AND Y = 74 else
"111111111111" when X = 230 AND Y = 74 else
"111111111111" when X = 231 AND Y = 74 else
"111111111111" when X = 232 AND Y = 74 else
"111111111111" when X = 233 AND Y = 74 else
"111111111111" when X = 234 AND Y = 74 else
"111111111111" when X = 235 AND Y = 74 else
"111111111111" when X = 236 AND Y = 74 else
"111111111111" when X = 237 AND Y = 74 else
"111111111111" when X = 238 AND Y = 74 else
"111111111111" when X = 239 AND Y = 74 else
"111111111111" when X = 240 AND Y = 74 else
"111111111111" when X = 241 AND Y = 74 else
"111111111111" when X = 242 AND Y = 74 else
"111111111111" when X = 243 AND Y = 74 else
"111111111111" when X = 244 AND Y = 74 else
"111111111111" when X = 245 AND Y = 74 else
"111111111111" when X = 246 AND Y = 74 else
"111111111111" when X = 247 AND Y = 74 else
"111111111111" when X = 248 AND Y = 74 else
"111111111111" when X = 249 AND Y = 74 else
"111111111111" when X = 250 AND Y = 74 else
"111111111111" when X = 251 AND Y = 74 else
"111111111111" when X = 252 AND Y = 74 else
"111111111111" when X = 253 AND Y = 74 else
"111111111111" when X = 254 AND Y = 74 else
"111111111111" when X = 255 AND Y = 74 else
"111111111111" when X = 256 AND Y = 74 else
"111111111111" when X = 257 AND Y = 74 else
"111111111111" when X = 258 AND Y = 74 else
"111111111111" when X = 259 AND Y = 74 else
"111111111111" when X = 260 AND Y = 74 else
"111111111111" when X = 261 AND Y = 74 else
"111111111111" when X = 262 AND Y = 74 else
"111111111111" when X = 263 AND Y = 74 else
"111111111111" when X = 264 AND Y = 74 else
"110111011111" when X = 265 AND Y = 74 else
"110111011111" when X = 266 AND Y = 74 else
"110111011111" when X = 267 AND Y = 74 else
"110111011111" when X = 268 AND Y = 74 else
"110111011111" when X = 269 AND Y = 74 else
"110111011111" when X = 270 AND Y = 74 else
"110111011111" when X = 271 AND Y = 74 else
"110111011111" when X = 272 AND Y = 74 else
"110111011111" when X = 273 AND Y = 74 else
"110111011111" when X = 274 AND Y = 74 else
"110111011111" when X = 275 AND Y = 74 else
"110111011111" when X = 276 AND Y = 74 else
"110111011111" when X = 277 AND Y = 74 else
"110111011111" when X = 278 AND Y = 74 else
"110111011111" when X = 279 AND Y = 74 else
"000000000000" when X = 280 AND Y = 74 else
"000000000000" when X = 281 AND Y = 74 else
"000000000000" when X = 282 AND Y = 74 else
"000000000000" when X = 283 AND Y = 74 else
"000000000000" when X = 284 AND Y = 74 else
"000000000000" when X = 285 AND Y = 74 else
"000000000000" when X = 286 AND Y = 74 else
"000000000000" when X = 287 AND Y = 74 else
"000000000000" when X = 288 AND Y = 74 else
"000000000000" when X = 289 AND Y = 74 else
"000000000000" when X = 290 AND Y = 74 else
"000000000000" when X = 291 AND Y = 74 else
"000000000000" when X = 292 AND Y = 74 else
"000000000000" when X = 293 AND Y = 74 else
"000000000000" when X = 294 AND Y = 74 else
"000000000000" when X = 295 AND Y = 74 else
"000000000000" when X = 296 AND Y = 74 else
"000000000000" when X = 297 AND Y = 74 else
"000000000000" when X = 298 AND Y = 74 else
"000000000000" when X = 299 AND Y = 74 else
"000000000000" when X = 300 AND Y = 74 else
"000000000000" when X = 301 AND Y = 74 else
"000000000000" when X = 302 AND Y = 74 else
"000000000000" when X = 303 AND Y = 74 else
"000000000000" when X = 304 AND Y = 74 else
"000000000000" when X = 305 AND Y = 74 else
"000000000000" when X = 306 AND Y = 74 else
"000000000000" when X = 307 AND Y = 74 else
"000000000000" when X = 308 AND Y = 74 else
"000000000000" when X = 309 AND Y = 74 else
"000000000000" when X = 310 AND Y = 74 else
"000000000000" when X = 311 AND Y = 74 else
"000000000000" when X = 312 AND Y = 74 else
"000000000000" when X = 313 AND Y = 74 else
"000000000000" when X = 314 AND Y = 74 else
"000000000000" when X = 315 AND Y = 74 else
"000000000000" when X = 316 AND Y = 74 else
"000000000000" when X = 317 AND Y = 74 else
"000000000000" when X = 318 AND Y = 74 else
"000000000000" when X = 319 AND Y = 74 else
"000000000000" when X = 320 AND Y = 74 else
"000000000000" when X = 321 AND Y = 74 else
"000000000000" when X = 322 AND Y = 74 else
"000000000000" when X = 323 AND Y = 74 else
"000000000000" when X = 324 AND Y = 74 else
"100010011101" when X = 0 AND Y = 75 else
"100010011101" when X = 1 AND Y = 75 else
"100010011101" when X = 2 AND Y = 75 else
"100010011101" when X = 3 AND Y = 75 else
"100010011101" when X = 4 AND Y = 75 else
"100010011101" when X = 5 AND Y = 75 else
"100010011101" when X = 6 AND Y = 75 else
"100010011101" when X = 7 AND Y = 75 else
"100010011101" when X = 8 AND Y = 75 else
"100010011101" when X = 9 AND Y = 75 else
"100010011101" when X = 10 AND Y = 75 else
"100010011101" when X = 11 AND Y = 75 else
"100010011101" when X = 12 AND Y = 75 else
"100010011101" when X = 13 AND Y = 75 else
"100010011101" when X = 14 AND Y = 75 else
"100010011101" when X = 15 AND Y = 75 else
"100010011101" when X = 16 AND Y = 75 else
"100010011101" when X = 17 AND Y = 75 else
"100010011101" when X = 18 AND Y = 75 else
"100010011101" when X = 19 AND Y = 75 else
"100010011101" when X = 20 AND Y = 75 else
"100010011101" when X = 21 AND Y = 75 else
"100010011101" when X = 22 AND Y = 75 else
"100010011101" when X = 23 AND Y = 75 else
"100010011101" when X = 24 AND Y = 75 else
"100010011101" when X = 25 AND Y = 75 else
"100010011101" when X = 26 AND Y = 75 else
"100010011101" when X = 27 AND Y = 75 else
"100010011101" when X = 28 AND Y = 75 else
"100010011101" when X = 29 AND Y = 75 else
"110111011111" when X = 30 AND Y = 75 else
"110111011111" when X = 31 AND Y = 75 else
"110111011111" when X = 32 AND Y = 75 else
"110111011111" when X = 33 AND Y = 75 else
"110111011111" when X = 34 AND Y = 75 else
"110111011111" when X = 35 AND Y = 75 else
"110111011111" when X = 36 AND Y = 75 else
"110111011111" when X = 37 AND Y = 75 else
"110111011111" when X = 38 AND Y = 75 else
"110111011111" when X = 39 AND Y = 75 else
"110111011111" when X = 40 AND Y = 75 else
"110111011111" when X = 41 AND Y = 75 else
"110111011111" when X = 42 AND Y = 75 else
"110111011111" when X = 43 AND Y = 75 else
"110111011111" when X = 44 AND Y = 75 else
"110111011111" when X = 45 AND Y = 75 else
"110111011111" when X = 46 AND Y = 75 else
"110111011111" when X = 47 AND Y = 75 else
"110111011111" when X = 48 AND Y = 75 else
"110111011111" when X = 49 AND Y = 75 else
"110111011111" when X = 50 AND Y = 75 else
"110111011111" when X = 51 AND Y = 75 else
"110111011111" when X = 52 AND Y = 75 else
"110111011111" when X = 53 AND Y = 75 else
"110111011111" when X = 54 AND Y = 75 else
"110111011111" when X = 55 AND Y = 75 else
"110111011111" when X = 56 AND Y = 75 else
"110111011111" when X = 57 AND Y = 75 else
"110111011111" when X = 58 AND Y = 75 else
"110111011111" when X = 59 AND Y = 75 else
"110111011111" when X = 60 AND Y = 75 else
"110111011111" when X = 61 AND Y = 75 else
"110111011111" when X = 62 AND Y = 75 else
"110111011111" when X = 63 AND Y = 75 else
"110111011111" when X = 64 AND Y = 75 else
"110111011111" when X = 65 AND Y = 75 else
"110111011111" when X = 66 AND Y = 75 else
"110111011111" when X = 67 AND Y = 75 else
"110111011111" when X = 68 AND Y = 75 else
"110111011111" when X = 69 AND Y = 75 else
"110111011111" when X = 70 AND Y = 75 else
"110111011111" when X = 71 AND Y = 75 else
"110111011111" when X = 72 AND Y = 75 else
"110111011111" when X = 73 AND Y = 75 else
"110111011111" when X = 74 AND Y = 75 else
"110111011111" when X = 75 AND Y = 75 else
"110111011111" when X = 76 AND Y = 75 else
"110111011111" when X = 77 AND Y = 75 else
"110111011111" when X = 78 AND Y = 75 else
"110111011111" when X = 79 AND Y = 75 else
"110111011111" when X = 80 AND Y = 75 else
"110111011111" when X = 81 AND Y = 75 else
"110111011111" when X = 82 AND Y = 75 else
"110111011111" when X = 83 AND Y = 75 else
"110111011111" when X = 84 AND Y = 75 else
"110111011111" when X = 85 AND Y = 75 else
"110111011111" when X = 86 AND Y = 75 else
"110111011111" when X = 87 AND Y = 75 else
"110111011111" when X = 88 AND Y = 75 else
"110111011111" when X = 89 AND Y = 75 else
"110111011111" when X = 90 AND Y = 75 else
"110111011111" when X = 91 AND Y = 75 else
"110111011111" when X = 92 AND Y = 75 else
"110111011111" when X = 93 AND Y = 75 else
"110111011111" when X = 94 AND Y = 75 else
"110111011111" when X = 95 AND Y = 75 else
"110111011111" when X = 96 AND Y = 75 else
"110111011111" when X = 97 AND Y = 75 else
"110111011111" when X = 98 AND Y = 75 else
"110111011111" when X = 99 AND Y = 75 else
"110111011111" when X = 100 AND Y = 75 else
"110111011111" when X = 101 AND Y = 75 else
"110111011111" when X = 102 AND Y = 75 else
"110111011111" when X = 103 AND Y = 75 else
"110111011111" when X = 104 AND Y = 75 else
"110111011111" when X = 105 AND Y = 75 else
"110111011111" when X = 106 AND Y = 75 else
"110111011111" when X = 107 AND Y = 75 else
"110111011111" when X = 108 AND Y = 75 else
"110111011111" when X = 109 AND Y = 75 else
"111111111111" when X = 110 AND Y = 75 else
"111111111111" when X = 111 AND Y = 75 else
"111111111111" when X = 112 AND Y = 75 else
"111111111111" when X = 113 AND Y = 75 else
"111111111111" when X = 114 AND Y = 75 else
"111111111111" when X = 115 AND Y = 75 else
"111111111111" when X = 116 AND Y = 75 else
"111111111111" when X = 117 AND Y = 75 else
"111111111111" when X = 118 AND Y = 75 else
"111111111111" when X = 119 AND Y = 75 else
"111111111111" when X = 120 AND Y = 75 else
"111111111111" when X = 121 AND Y = 75 else
"111111111111" when X = 122 AND Y = 75 else
"111111111111" when X = 123 AND Y = 75 else
"111111111111" when X = 124 AND Y = 75 else
"111111111111" when X = 125 AND Y = 75 else
"111111111111" when X = 126 AND Y = 75 else
"111111111111" when X = 127 AND Y = 75 else
"111111111111" when X = 128 AND Y = 75 else
"111111111111" when X = 129 AND Y = 75 else
"111111111111" when X = 130 AND Y = 75 else
"111111111111" when X = 131 AND Y = 75 else
"111111111111" when X = 132 AND Y = 75 else
"111111111111" when X = 133 AND Y = 75 else
"111111111111" when X = 134 AND Y = 75 else
"111111111111" when X = 135 AND Y = 75 else
"111111111111" when X = 136 AND Y = 75 else
"111111111111" when X = 137 AND Y = 75 else
"111111111111" when X = 138 AND Y = 75 else
"111111111111" when X = 139 AND Y = 75 else
"111111111111" when X = 140 AND Y = 75 else
"111111111111" when X = 141 AND Y = 75 else
"111111111111" when X = 142 AND Y = 75 else
"111111111111" when X = 143 AND Y = 75 else
"111111111111" when X = 144 AND Y = 75 else
"111111111111" when X = 145 AND Y = 75 else
"111111111111" when X = 146 AND Y = 75 else
"111111111111" when X = 147 AND Y = 75 else
"111111111111" when X = 148 AND Y = 75 else
"111111111111" when X = 149 AND Y = 75 else
"111111111111" when X = 150 AND Y = 75 else
"111111111111" when X = 151 AND Y = 75 else
"111111111111" when X = 152 AND Y = 75 else
"111111111111" when X = 153 AND Y = 75 else
"111111111111" when X = 154 AND Y = 75 else
"111111111111" when X = 155 AND Y = 75 else
"111111111111" when X = 156 AND Y = 75 else
"111111111111" when X = 157 AND Y = 75 else
"111111111111" when X = 158 AND Y = 75 else
"111111111111" when X = 159 AND Y = 75 else
"111111111111" when X = 160 AND Y = 75 else
"111111111111" when X = 161 AND Y = 75 else
"111111111111" when X = 162 AND Y = 75 else
"111111111111" when X = 163 AND Y = 75 else
"111111111111" when X = 164 AND Y = 75 else
"111111111111" when X = 165 AND Y = 75 else
"111111111111" when X = 166 AND Y = 75 else
"111111111111" when X = 167 AND Y = 75 else
"111111111111" when X = 168 AND Y = 75 else
"111111111111" when X = 169 AND Y = 75 else
"111111111111" when X = 170 AND Y = 75 else
"111111111111" when X = 171 AND Y = 75 else
"111111111111" when X = 172 AND Y = 75 else
"111111111111" when X = 173 AND Y = 75 else
"111111111111" when X = 174 AND Y = 75 else
"111111111111" when X = 175 AND Y = 75 else
"111111111111" when X = 176 AND Y = 75 else
"111111111111" when X = 177 AND Y = 75 else
"111111111111" when X = 178 AND Y = 75 else
"111111111111" when X = 179 AND Y = 75 else
"111111111111" when X = 180 AND Y = 75 else
"111111111111" when X = 181 AND Y = 75 else
"111111111111" when X = 182 AND Y = 75 else
"111111111111" when X = 183 AND Y = 75 else
"111111111111" when X = 184 AND Y = 75 else
"111111111111" when X = 185 AND Y = 75 else
"111111111111" when X = 186 AND Y = 75 else
"111111111111" when X = 187 AND Y = 75 else
"111111111111" when X = 188 AND Y = 75 else
"111111111111" when X = 189 AND Y = 75 else
"111111111111" when X = 190 AND Y = 75 else
"111111111111" when X = 191 AND Y = 75 else
"111111111111" when X = 192 AND Y = 75 else
"111111111111" when X = 193 AND Y = 75 else
"111111111111" when X = 194 AND Y = 75 else
"111111111111" when X = 195 AND Y = 75 else
"111111111111" when X = 196 AND Y = 75 else
"111111111111" when X = 197 AND Y = 75 else
"111111111111" when X = 198 AND Y = 75 else
"111111111111" when X = 199 AND Y = 75 else
"111111111111" when X = 200 AND Y = 75 else
"111111111111" when X = 201 AND Y = 75 else
"111111111111" when X = 202 AND Y = 75 else
"111111111111" when X = 203 AND Y = 75 else
"111111111111" when X = 204 AND Y = 75 else
"111111111111" when X = 205 AND Y = 75 else
"111111111111" when X = 206 AND Y = 75 else
"111111111111" when X = 207 AND Y = 75 else
"111111111111" when X = 208 AND Y = 75 else
"111111111111" when X = 209 AND Y = 75 else
"111111111111" when X = 210 AND Y = 75 else
"111111111111" when X = 211 AND Y = 75 else
"111111111111" when X = 212 AND Y = 75 else
"111111111111" when X = 213 AND Y = 75 else
"111111111111" when X = 214 AND Y = 75 else
"111111111111" when X = 215 AND Y = 75 else
"111111111111" when X = 216 AND Y = 75 else
"111111111111" when X = 217 AND Y = 75 else
"111111111111" when X = 218 AND Y = 75 else
"111111111111" when X = 219 AND Y = 75 else
"111111111111" when X = 220 AND Y = 75 else
"111111111111" when X = 221 AND Y = 75 else
"111111111111" when X = 222 AND Y = 75 else
"111111111111" when X = 223 AND Y = 75 else
"111111111111" when X = 224 AND Y = 75 else
"111111111111" when X = 225 AND Y = 75 else
"111111111111" when X = 226 AND Y = 75 else
"111111111111" when X = 227 AND Y = 75 else
"111111111111" when X = 228 AND Y = 75 else
"111111111111" when X = 229 AND Y = 75 else
"111111111111" when X = 230 AND Y = 75 else
"111111111111" when X = 231 AND Y = 75 else
"111111111111" when X = 232 AND Y = 75 else
"111111111111" when X = 233 AND Y = 75 else
"111111111111" when X = 234 AND Y = 75 else
"111111111111" when X = 235 AND Y = 75 else
"111111111111" when X = 236 AND Y = 75 else
"111111111111" when X = 237 AND Y = 75 else
"111111111111" when X = 238 AND Y = 75 else
"111111111111" when X = 239 AND Y = 75 else
"111111111111" when X = 240 AND Y = 75 else
"111111111111" when X = 241 AND Y = 75 else
"111111111111" when X = 242 AND Y = 75 else
"111111111111" when X = 243 AND Y = 75 else
"111111111111" when X = 244 AND Y = 75 else
"111111111111" when X = 245 AND Y = 75 else
"111111111111" when X = 246 AND Y = 75 else
"111111111111" when X = 247 AND Y = 75 else
"111111111111" when X = 248 AND Y = 75 else
"111111111111" when X = 249 AND Y = 75 else
"111111111111" when X = 250 AND Y = 75 else
"111111111111" when X = 251 AND Y = 75 else
"111111111111" when X = 252 AND Y = 75 else
"111111111111" when X = 253 AND Y = 75 else
"111111111111" when X = 254 AND Y = 75 else
"111111111111" when X = 255 AND Y = 75 else
"111111111111" when X = 256 AND Y = 75 else
"111111111111" when X = 257 AND Y = 75 else
"111111111111" when X = 258 AND Y = 75 else
"111111111111" when X = 259 AND Y = 75 else
"111111111111" when X = 260 AND Y = 75 else
"111111111111" when X = 261 AND Y = 75 else
"111111111111" when X = 262 AND Y = 75 else
"111111111111" when X = 263 AND Y = 75 else
"111111111111" when X = 264 AND Y = 75 else
"110111011111" when X = 265 AND Y = 75 else
"110111011111" when X = 266 AND Y = 75 else
"110111011111" when X = 267 AND Y = 75 else
"110111011111" when X = 268 AND Y = 75 else
"110111011111" when X = 269 AND Y = 75 else
"110111011111" when X = 270 AND Y = 75 else
"110111011111" when X = 271 AND Y = 75 else
"110111011111" when X = 272 AND Y = 75 else
"110111011111" when X = 273 AND Y = 75 else
"110111011111" when X = 274 AND Y = 75 else
"110111011111" when X = 275 AND Y = 75 else
"110111011111" when X = 276 AND Y = 75 else
"110111011111" when X = 277 AND Y = 75 else
"110111011111" when X = 278 AND Y = 75 else
"110111011111" when X = 279 AND Y = 75 else
"000000000000" when X = 280 AND Y = 75 else
"000000000000" when X = 281 AND Y = 75 else
"000000000000" when X = 282 AND Y = 75 else
"000000000000" when X = 283 AND Y = 75 else
"000000000000" when X = 284 AND Y = 75 else
"000000000000" when X = 285 AND Y = 75 else
"000000000000" when X = 286 AND Y = 75 else
"000000000000" when X = 287 AND Y = 75 else
"000000000000" when X = 288 AND Y = 75 else
"000000000000" when X = 289 AND Y = 75 else
"000000000000" when X = 290 AND Y = 75 else
"000000000000" when X = 291 AND Y = 75 else
"000000000000" when X = 292 AND Y = 75 else
"000000000000" when X = 293 AND Y = 75 else
"000000000000" when X = 294 AND Y = 75 else
"000000000000" when X = 295 AND Y = 75 else
"000000000000" when X = 296 AND Y = 75 else
"000000000000" when X = 297 AND Y = 75 else
"000000000000" when X = 298 AND Y = 75 else
"000000000000" when X = 299 AND Y = 75 else
"000000000000" when X = 300 AND Y = 75 else
"000000000000" when X = 301 AND Y = 75 else
"000000000000" when X = 302 AND Y = 75 else
"000000000000" when X = 303 AND Y = 75 else
"000000000000" when X = 304 AND Y = 75 else
"000000000000" when X = 305 AND Y = 75 else
"000000000000" when X = 306 AND Y = 75 else
"000000000000" when X = 307 AND Y = 75 else
"000000000000" when X = 308 AND Y = 75 else
"000000000000" when X = 309 AND Y = 75 else
"000000000000" when X = 310 AND Y = 75 else
"000000000000" when X = 311 AND Y = 75 else
"000000000000" when X = 312 AND Y = 75 else
"000000000000" when X = 313 AND Y = 75 else
"000000000000" when X = 314 AND Y = 75 else
"000000000000" when X = 315 AND Y = 75 else
"000000000000" when X = 316 AND Y = 75 else
"000000000000" when X = 317 AND Y = 75 else
"000000000000" when X = 318 AND Y = 75 else
"000000000000" when X = 319 AND Y = 75 else
"000000000000" when X = 320 AND Y = 75 else
"000000000000" when X = 321 AND Y = 75 else
"000000000000" when X = 322 AND Y = 75 else
"000000000000" when X = 323 AND Y = 75 else
"000000000000" when X = 324 AND Y = 75 else
"100010011101" when X = 0 AND Y = 76 else
"100010011101" when X = 1 AND Y = 76 else
"100010011101" when X = 2 AND Y = 76 else
"100010011101" when X = 3 AND Y = 76 else
"100010011101" when X = 4 AND Y = 76 else
"100010011101" when X = 5 AND Y = 76 else
"100010011101" when X = 6 AND Y = 76 else
"100010011101" when X = 7 AND Y = 76 else
"100010011101" when X = 8 AND Y = 76 else
"100010011101" when X = 9 AND Y = 76 else
"100010011101" when X = 10 AND Y = 76 else
"100010011101" when X = 11 AND Y = 76 else
"100010011101" when X = 12 AND Y = 76 else
"100010011101" when X = 13 AND Y = 76 else
"100010011101" when X = 14 AND Y = 76 else
"100010011101" when X = 15 AND Y = 76 else
"100010011101" when X = 16 AND Y = 76 else
"100010011101" when X = 17 AND Y = 76 else
"100010011101" when X = 18 AND Y = 76 else
"100010011101" when X = 19 AND Y = 76 else
"100010011101" when X = 20 AND Y = 76 else
"100010011101" when X = 21 AND Y = 76 else
"100010011101" when X = 22 AND Y = 76 else
"100010011101" when X = 23 AND Y = 76 else
"100010011101" when X = 24 AND Y = 76 else
"100010011101" when X = 25 AND Y = 76 else
"100010011101" when X = 26 AND Y = 76 else
"100010011101" when X = 27 AND Y = 76 else
"100010011101" when X = 28 AND Y = 76 else
"100010011101" when X = 29 AND Y = 76 else
"110111011111" when X = 30 AND Y = 76 else
"110111011111" when X = 31 AND Y = 76 else
"110111011111" when X = 32 AND Y = 76 else
"110111011111" when X = 33 AND Y = 76 else
"110111011111" when X = 34 AND Y = 76 else
"110111011111" when X = 35 AND Y = 76 else
"110111011111" when X = 36 AND Y = 76 else
"110111011111" when X = 37 AND Y = 76 else
"110111011111" when X = 38 AND Y = 76 else
"110111011111" when X = 39 AND Y = 76 else
"110111011111" when X = 40 AND Y = 76 else
"110111011111" when X = 41 AND Y = 76 else
"110111011111" when X = 42 AND Y = 76 else
"110111011111" when X = 43 AND Y = 76 else
"110111011111" when X = 44 AND Y = 76 else
"110111011111" when X = 45 AND Y = 76 else
"110111011111" when X = 46 AND Y = 76 else
"110111011111" when X = 47 AND Y = 76 else
"110111011111" when X = 48 AND Y = 76 else
"110111011111" when X = 49 AND Y = 76 else
"110111011111" when X = 50 AND Y = 76 else
"110111011111" when X = 51 AND Y = 76 else
"110111011111" when X = 52 AND Y = 76 else
"110111011111" when X = 53 AND Y = 76 else
"110111011111" when X = 54 AND Y = 76 else
"110111011111" when X = 55 AND Y = 76 else
"110111011111" when X = 56 AND Y = 76 else
"110111011111" when X = 57 AND Y = 76 else
"110111011111" when X = 58 AND Y = 76 else
"110111011111" when X = 59 AND Y = 76 else
"110111011111" when X = 60 AND Y = 76 else
"110111011111" when X = 61 AND Y = 76 else
"110111011111" when X = 62 AND Y = 76 else
"110111011111" when X = 63 AND Y = 76 else
"110111011111" when X = 64 AND Y = 76 else
"110111011111" when X = 65 AND Y = 76 else
"110111011111" when X = 66 AND Y = 76 else
"110111011111" when X = 67 AND Y = 76 else
"110111011111" when X = 68 AND Y = 76 else
"110111011111" when X = 69 AND Y = 76 else
"110111011111" when X = 70 AND Y = 76 else
"110111011111" when X = 71 AND Y = 76 else
"110111011111" when X = 72 AND Y = 76 else
"110111011111" when X = 73 AND Y = 76 else
"110111011111" when X = 74 AND Y = 76 else
"110111011111" when X = 75 AND Y = 76 else
"110111011111" when X = 76 AND Y = 76 else
"110111011111" when X = 77 AND Y = 76 else
"110111011111" when X = 78 AND Y = 76 else
"110111011111" when X = 79 AND Y = 76 else
"110111011111" when X = 80 AND Y = 76 else
"110111011111" when X = 81 AND Y = 76 else
"110111011111" when X = 82 AND Y = 76 else
"110111011111" when X = 83 AND Y = 76 else
"110111011111" when X = 84 AND Y = 76 else
"110111011111" when X = 85 AND Y = 76 else
"110111011111" when X = 86 AND Y = 76 else
"110111011111" when X = 87 AND Y = 76 else
"110111011111" when X = 88 AND Y = 76 else
"110111011111" when X = 89 AND Y = 76 else
"110111011111" when X = 90 AND Y = 76 else
"110111011111" when X = 91 AND Y = 76 else
"110111011111" when X = 92 AND Y = 76 else
"110111011111" when X = 93 AND Y = 76 else
"110111011111" when X = 94 AND Y = 76 else
"110111011111" when X = 95 AND Y = 76 else
"110111011111" when X = 96 AND Y = 76 else
"110111011111" when X = 97 AND Y = 76 else
"110111011111" when X = 98 AND Y = 76 else
"110111011111" when X = 99 AND Y = 76 else
"110111011111" when X = 100 AND Y = 76 else
"110111011111" when X = 101 AND Y = 76 else
"110111011111" when X = 102 AND Y = 76 else
"110111011111" when X = 103 AND Y = 76 else
"110111011111" when X = 104 AND Y = 76 else
"110111011111" when X = 105 AND Y = 76 else
"110111011111" when X = 106 AND Y = 76 else
"110111011111" when X = 107 AND Y = 76 else
"110111011111" when X = 108 AND Y = 76 else
"110111011111" when X = 109 AND Y = 76 else
"111111111111" when X = 110 AND Y = 76 else
"111111111111" when X = 111 AND Y = 76 else
"111111111111" when X = 112 AND Y = 76 else
"111111111111" when X = 113 AND Y = 76 else
"111111111111" when X = 114 AND Y = 76 else
"111111111111" when X = 115 AND Y = 76 else
"111111111111" when X = 116 AND Y = 76 else
"111111111111" when X = 117 AND Y = 76 else
"111111111111" when X = 118 AND Y = 76 else
"111111111111" when X = 119 AND Y = 76 else
"111111111111" when X = 120 AND Y = 76 else
"111111111111" when X = 121 AND Y = 76 else
"111111111111" when X = 122 AND Y = 76 else
"111111111111" when X = 123 AND Y = 76 else
"111111111111" when X = 124 AND Y = 76 else
"111111111111" when X = 125 AND Y = 76 else
"111111111111" when X = 126 AND Y = 76 else
"111111111111" when X = 127 AND Y = 76 else
"111111111111" when X = 128 AND Y = 76 else
"111111111111" when X = 129 AND Y = 76 else
"111111111111" when X = 130 AND Y = 76 else
"111111111111" when X = 131 AND Y = 76 else
"111111111111" when X = 132 AND Y = 76 else
"111111111111" when X = 133 AND Y = 76 else
"111111111111" when X = 134 AND Y = 76 else
"111111111111" when X = 135 AND Y = 76 else
"111111111111" when X = 136 AND Y = 76 else
"111111111111" when X = 137 AND Y = 76 else
"111111111111" when X = 138 AND Y = 76 else
"111111111111" when X = 139 AND Y = 76 else
"111111111111" when X = 140 AND Y = 76 else
"111111111111" when X = 141 AND Y = 76 else
"111111111111" when X = 142 AND Y = 76 else
"111111111111" when X = 143 AND Y = 76 else
"111111111111" when X = 144 AND Y = 76 else
"111111111111" when X = 145 AND Y = 76 else
"111111111111" when X = 146 AND Y = 76 else
"111111111111" when X = 147 AND Y = 76 else
"111111111111" when X = 148 AND Y = 76 else
"111111111111" when X = 149 AND Y = 76 else
"111111111111" when X = 150 AND Y = 76 else
"111111111111" when X = 151 AND Y = 76 else
"111111111111" when X = 152 AND Y = 76 else
"111111111111" when X = 153 AND Y = 76 else
"111111111111" when X = 154 AND Y = 76 else
"111111111111" when X = 155 AND Y = 76 else
"111111111111" when X = 156 AND Y = 76 else
"111111111111" when X = 157 AND Y = 76 else
"111111111111" when X = 158 AND Y = 76 else
"111111111111" when X = 159 AND Y = 76 else
"111111111111" when X = 160 AND Y = 76 else
"111111111111" when X = 161 AND Y = 76 else
"111111111111" when X = 162 AND Y = 76 else
"111111111111" when X = 163 AND Y = 76 else
"111111111111" when X = 164 AND Y = 76 else
"111111111111" when X = 165 AND Y = 76 else
"111111111111" when X = 166 AND Y = 76 else
"111111111111" when X = 167 AND Y = 76 else
"111111111111" when X = 168 AND Y = 76 else
"111111111111" when X = 169 AND Y = 76 else
"111111111111" when X = 170 AND Y = 76 else
"111111111111" when X = 171 AND Y = 76 else
"111111111111" when X = 172 AND Y = 76 else
"111111111111" when X = 173 AND Y = 76 else
"111111111111" when X = 174 AND Y = 76 else
"111111111111" when X = 175 AND Y = 76 else
"111111111111" when X = 176 AND Y = 76 else
"111111111111" when X = 177 AND Y = 76 else
"111111111111" when X = 178 AND Y = 76 else
"111111111111" when X = 179 AND Y = 76 else
"111111111111" when X = 180 AND Y = 76 else
"111111111111" when X = 181 AND Y = 76 else
"111111111111" when X = 182 AND Y = 76 else
"111111111111" when X = 183 AND Y = 76 else
"111111111111" when X = 184 AND Y = 76 else
"111111111111" when X = 185 AND Y = 76 else
"111111111111" when X = 186 AND Y = 76 else
"111111111111" when X = 187 AND Y = 76 else
"111111111111" when X = 188 AND Y = 76 else
"111111111111" when X = 189 AND Y = 76 else
"111111111111" when X = 190 AND Y = 76 else
"111111111111" when X = 191 AND Y = 76 else
"111111111111" when X = 192 AND Y = 76 else
"111111111111" when X = 193 AND Y = 76 else
"111111111111" when X = 194 AND Y = 76 else
"111111111111" when X = 195 AND Y = 76 else
"111111111111" when X = 196 AND Y = 76 else
"111111111111" when X = 197 AND Y = 76 else
"111111111111" when X = 198 AND Y = 76 else
"111111111111" when X = 199 AND Y = 76 else
"111111111111" when X = 200 AND Y = 76 else
"111111111111" when X = 201 AND Y = 76 else
"111111111111" when X = 202 AND Y = 76 else
"111111111111" when X = 203 AND Y = 76 else
"111111111111" when X = 204 AND Y = 76 else
"111111111111" when X = 205 AND Y = 76 else
"111111111111" when X = 206 AND Y = 76 else
"111111111111" when X = 207 AND Y = 76 else
"111111111111" when X = 208 AND Y = 76 else
"111111111111" when X = 209 AND Y = 76 else
"111111111111" when X = 210 AND Y = 76 else
"111111111111" when X = 211 AND Y = 76 else
"111111111111" when X = 212 AND Y = 76 else
"111111111111" when X = 213 AND Y = 76 else
"111111111111" when X = 214 AND Y = 76 else
"111111111111" when X = 215 AND Y = 76 else
"111111111111" when X = 216 AND Y = 76 else
"111111111111" when X = 217 AND Y = 76 else
"111111111111" when X = 218 AND Y = 76 else
"111111111111" when X = 219 AND Y = 76 else
"111111111111" when X = 220 AND Y = 76 else
"111111111111" when X = 221 AND Y = 76 else
"111111111111" when X = 222 AND Y = 76 else
"111111111111" when X = 223 AND Y = 76 else
"111111111111" when X = 224 AND Y = 76 else
"111111111111" when X = 225 AND Y = 76 else
"111111111111" when X = 226 AND Y = 76 else
"111111111111" when X = 227 AND Y = 76 else
"111111111111" when X = 228 AND Y = 76 else
"111111111111" when X = 229 AND Y = 76 else
"111111111111" when X = 230 AND Y = 76 else
"111111111111" when X = 231 AND Y = 76 else
"111111111111" when X = 232 AND Y = 76 else
"111111111111" when X = 233 AND Y = 76 else
"111111111111" when X = 234 AND Y = 76 else
"111111111111" when X = 235 AND Y = 76 else
"111111111111" when X = 236 AND Y = 76 else
"111111111111" when X = 237 AND Y = 76 else
"111111111111" when X = 238 AND Y = 76 else
"111111111111" when X = 239 AND Y = 76 else
"111111111111" when X = 240 AND Y = 76 else
"111111111111" when X = 241 AND Y = 76 else
"111111111111" when X = 242 AND Y = 76 else
"111111111111" when X = 243 AND Y = 76 else
"111111111111" when X = 244 AND Y = 76 else
"111111111111" when X = 245 AND Y = 76 else
"111111111111" when X = 246 AND Y = 76 else
"111111111111" when X = 247 AND Y = 76 else
"111111111111" when X = 248 AND Y = 76 else
"111111111111" when X = 249 AND Y = 76 else
"111111111111" when X = 250 AND Y = 76 else
"111111111111" when X = 251 AND Y = 76 else
"111111111111" when X = 252 AND Y = 76 else
"111111111111" when X = 253 AND Y = 76 else
"111111111111" when X = 254 AND Y = 76 else
"111111111111" when X = 255 AND Y = 76 else
"111111111111" when X = 256 AND Y = 76 else
"111111111111" when X = 257 AND Y = 76 else
"111111111111" when X = 258 AND Y = 76 else
"111111111111" when X = 259 AND Y = 76 else
"111111111111" when X = 260 AND Y = 76 else
"111111111111" when X = 261 AND Y = 76 else
"111111111111" when X = 262 AND Y = 76 else
"111111111111" when X = 263 AND Y = 76 else
"111111111111" when X = 264 AND Y = 76 else
"110111011111" when X = 265 AND Y = 76 else
"110111011111" when X = 266 AND Y = 76 else
"110111011111" when X = 267 AND Y = 76 else
"110111011111" when X = 268 AND Y = 76 else
"110111011111" when X = 269 AND Y = 76 else
"110111011111" when X = 270 AND Y = 76 else
"110111011111" when X = 271 AND Y = 76 else
"110111011111" when X = 272 AND Y = 76 else
"110111011111" when X = 273 AND Y = 76 else
"110111011111" when X = 274 AND Y = 76 else
"110111011111" when X = 275 AND Y = 76 else
"110111011111" when X = 276 AND Y = 76 else
"110111011111" when X = 277 AND Y = 76 else
"110111011111" when X = 278 AND Y = 76 else
"110111011111" when X = 279 AND Y = 76 else
"000000000000" when X = 280 AND Y = 76 else
"000000000000" when X = 281 AND Y = 76 else
"000000000000" when X = 282 AND Y = 76 else
"000000000000" when X = 283 AND Y = 76 else
"000000000000" when X = 284 AND Y = 76 else
"000000000000" when X = 285 AND Y = 76 else
"000000000000" when X = 286 AND Y = 76 else
"000000000000" when X = 287 AND Y = 76 else
"000000000000" when X = 288 AND Y = 76 else
"000000000000" when X = 289 AND Y = 76 else
"000000000000" when X = 290 AND Y = 76 else
"000000000000" when X = 291 AND Y = 76 else
"000000000000" when X = 292 AND Y = 76 else
"000000000000" when X = 293 AND Y = 76 else
"000000000000" when X = 294 AND Y = 76 else
"000000000000" when X = 295 AND Y = 76 else
"000000000000" when X = 296 AND Y = 76 else
"000000000000" when X = 297 AND Y = 76 else
"000000000000" when X = 298 AND Y = 76 else
"000000000000" when X = 299 AND Y = 76 else
"000000000000" when X = 300 AND Y = 76 else
"000000000000" when X = 301 AND Y = 76 else
"000000000000" when X = 302 AND Y = 76 else
"000000000000" when X = 303 AND Y = 76 else
"000000000000" when X = 304 AND Y = 76 else
"000000000000" when X = 305 AND Y = 76 else
"000000000000" when X = 306 AND Y = 76 else
"000000000000" when X = 307 AND Y = 76 else
"000000000000" when X = 308 AND Y = 76 else
"000000000000" when X = 309 AND Y = 76 else
"000000000000" when X = 310 AND Y = 76 else
"000000000000" when X = 311 AND Y = 76 else
"000000000000" when X = 312 AND Y = 76 else
"000000000000" when X = 313 AND Y = 76 else
"000000000000" when X = 314 AND Y = 76 else
"000000000000" when X = 315 AND Y = 76 else
"000000000000" when X = 316 AND Y = 76 else
"000000000000" when X = 317 AND Y = 76 else
"000000000000" when X = 318 AND Y = 76 else
"000000000000" when X = 319 AND Y = 76 else
"000000000000" when X = 320 AND Y = 76 else
"000000000000" when X = 321 AND Y = 76 else
"000000000000" when X = 322 AND Y = 76 else
"000000000000" when X = 323 AND Y = 76 else
"000000000000" when X = 324 AND Y = 76 else
"100010011101" when X = 0 AND Y = 77 else
"100010011101" when X = 1 AND Y = 77 else
"100010011101" when X = 2 AND Y = 77 else
"100010011101" when X = 3 AND Y = 77 else
"100010011101" when X = 4 AND Y = 77 else
"100010011101" when X = 5 AND Y = 77 else
"100010011101" when X = 6 AND Y = 77 else
"100010011101" when X = 7 AND Y = 77 else
"100010011101" when X = 8 AND Y = 77 else
"100010011101" when X = 9 AND Y = 77 else
"100010011101" when X = 10 AND Y = 77 else
"100010011101" when X = 11 AND Y = 77 else
"100010011101" when X = 12 AND Y = 77 else
"100010011101" when X = 13 AND Y = 77 else
"100010011101" when X = 14 AND Y = 77 else
"100010011101" when X = 15 AND Y = 77 else
"100010011101" when X = 16 AND Y = 77 else
"100010011101" when X = 17 AND Y = 77 else
"100010011101" when X = 18 AND Y = 77 else
"100010011101" when X = 19 AND Y = 77 else
"100010011101" when X = 20 AND Y = 77 else
"100010011101" when X = 21 AND Y = 77 else
"100010011101" when X = 22 AND Y = 77 else
"100010011101" when X = 23 AND Y = 77 else
"100010011101" when X = 24 AND Y = 77 else
"100010011101" when X = 25 AND Y = 77 else
"100010011101" when X = 26 AND Y = 77 else
"100010011101" when X = 27 AND Y = 77 else
"100010011101" when X = 28 AND Y = 77 else
"100010011101" when X = 29 AND Y = 77 else
"110111011111" when X = 30 AND Y = 77 else
"110111011111" when X = 31 AND Y = 77 else
"110111011111" when X = 32 AND Y = 77 else
"110111011111" when X = 33 AND Y = 77 else
"110111011111" when X = 34 AND Y = 77 else
"110111011111" when X = 35 AND Y = 77 else
"110111011111" when X = 36 AND Y = 77 else
"110111011111" when X = 37 AND Y = 77 else
"110111011111" when X = 38 AND Y = 77 else
"110111011111" when X = 39 AND Y = 77 else
"110111011111" when X = 40 AND Y = 77 else
"110111011111" when X = 41 AND Y = 77 else
"110111011111" when X = 42 AND Y = 77 else
"110111011111" when X = 43 AND Y = 77 else
"110111011111" when X = 44 AND Y = 77 else
"110111011111" when X = 45 AND Y = 77 else
"110111011111" when X = 46 AND Y = 77 else
"110111011111" when X = 47 AND Y = 77 else
"110111011111" when X = 48 AND Y = 77 else
"110111011111" when X = 49 AND Y = 77 else
"110111011111" when X = 50 AND Y = 77 else
"110111011111" when X = 51 AND Y = 77 else
"110111011111" when X = 52 AND Y = 77 else
"110111011111" when X = 53 AND Y = 77 else
"110111011111" when X = 54 AND Y = 77 else
"110111011111" when X = 55 AND Y = 77 else
"110111011111" when X = 56 AND Y = 77 else
"110111011111" when X = 57 AND Y = 77 else
"110111011111" when X = 58 AND Y = 77 else
"110111011111" when X = 59 AND Y = 77 else
"110111011111" when X = 60 AND Y = 77 else
"110111011111" when X = 61 AND Y = 77 else
"110111011111" when X = 62 AND Y = 77 else
"110111011111" when X = 63 AND Y = 77 else
"110111011111" when X = 64 AND Y = 77 else
"110111011111" when X = 65 AND Y = 77 else
"110111011111" when X = 66 AND Y = 77 else
"110111011111" when X = 67 AND Y = 77 else
"110111011111" when X = 68 AND Y = 77 else
"110111011111" when X = 69 AND Y = 77 else
"110111011111" when X = 70 AND Y = 77 else
"110111011111" when X = 71 AND Y = 77 else
"110111011111" when X = 72 AND Y = 77 else
"110111011111" when X = 73 AND Y = 77 else
"110111011111" when X = 74 AND Y = 77 else
"110111011111" when X = 75 AND Y = 77 else
"110111011111" when X = 76 AND Y = 77 else
"110111011111" when X = 77 AND Y = 77 else
"110111011111" when X = 78 AND Y = 77 else
"110111011111" when X = 79 AND Y = 77 else
"110111011111" when X = 80 AND Y = 77 else
"110111011111" when X = 81 AND Y = 77 else
"110111011111" when X = 82 AND Y = 77 else
"110111011111" when X = 83 AND Y = 77 else
"110111011111" when X = 84 AND Y = 77 else
"110111011111" when X = 85 AND Y = 77 else
"110111011111" when X = 86 AND Y = 77 else
"110111011111" when X = 87 AND Y = 77 else
"110111011111" when X = 88 AND Y = 77 else
"110111011111" when X = 89 AND Y = 77 else
"110111011111" when X = 90 AND Y = 77 else
"110111011111" when X = 91 AND Y = 77 else
"110111011111" when X = 92 AND Y = 77 else
"110111011111" when X = 93 AND Y = 77 else
"110111011111" when X = 94 AND Y = 77 else
"110111011111" when X = 95 AND Y = 77 else
"110111011111" when X = 96 AND Y = 77 else
"110111011111" when X = 97 AND Y = 77 else
"110111011111" when X = 98 AND Y = 77 else
"110111011111" when X = 99 AND Y = 77 else
"110111011111" when X = 100 AND Y = 77 else
"110111011111" when X = 101 AND Y = 77 else
"110111011111" when X = 102 AND Y = 77 else
"110111011111" when X = 103 AND Y = 77 else
"110111011111" when X = 104 AND Y = 77 else
"110111011111" when X = 105 AND Y = 77 else
"110111011111" when X = 106 AND Y = 77 else
"110111011111" when X = 107 AND Y = 77 else
"110111011111" when X = 108 AND Y = 77 else
"110111011111" when X = 109 AND Y = 77 else
"111111111111" when X = 110 AND Y = 77 else
"111111111111" when X = 111 AND Y = 77 else
"111111111111" when X = 112 AND Y = 77 else
"111111111111" when X = 113 AND Y = 77 else
"111111111111" when X = 114 AND Y = 77 else
"111111111111" when X = 115 AND Y = 77 else
"111111111111" when X = 116 AND Y = 77 else
"111111111111" when X = 117 AND Y = 77 else
"111111111111" when X = 118 AND Y = 77 else
"111111111111" when X = 119 AND Y = 77 else
"111111111111" when X = 120 AND Y = 77 else
"111111111111" when X = 121 AND Y = 77 else
"111111111111" when X = 122 AND Y = 77 else
"111111111111" when X = 123 AND Y = 77 else
"111111111111" when X = 124 AND Y = 77 else
"111111111111" when X = 125 AND Y = 77 else
"111111111111" when X = 126 AND Y = 77 else
"111111111111" when X = 127 AND Y = 77 else
"111111111111" when X = 128 AND Y = 77 else
"111111111111" when X = 129 AND Y = 77 else
"111111111111" when X = 130 AND Y = 77 else
"111111111111" when X = 131 AND Y = 77 else
"111111111111" when X = 132 AND Y = 77 else
"111111111111" when X = 133 AND Y = 77 else
"111111111111" when X = 134 AND Y = 77 else
"111111111111" when X = 135 AND Y = 77 else
"111111111111" when X = 136 AND Y = 77 else
"111111111111" when X = 137 AND Y = 77 else
"111111111111" when X = 138 AND Y = 77 else
"111111111111" when X = 139 AND Y = 77 else
"111111111111" when X = 140 AND Y = 77 else
"111111111111" when X = 141 AND Y = 77 else
"111111111111" when X = 142 AND Y = 77 else
"111111111111" when X = 143 AND Y = 77 else
"111111111111" when X = 144 AND Y = 77 else
"111111111111" when X = 145 AND Y = 77 else
"111111111111" when X = 146 AND Y = 77 else
"111111111111" when X = 147 AND Y = 77 else
"111111111111" when X = 148 AND Y = 77 else
"111111111111" when X = 149 AND Y = 77 else
"111111111111" when X = 150 AND Y = 77 else
"111111111111" when X = 151 AND Y = 77 else
"111111111111" when X = 152 AND Y = 77 else
"111111111111" when X = 153 AND Y = 77 else
"111111111111" when X = 154 AND Y = 77 else
"111111111111" when X = 155 AND Y = 77 else
"111111111111" when X = 156 AND Y = 77 else
"111111111111" when X = 157 AND Y = 77 else
"111111111111" when X = 158 AND Y = 77 else
"111111111111" when X = 159 AND Y = 77 else
"111111111111" when X = 160 AND Y = 77 else
"111111111111" when X = 161 AND Y = 77 else
"111111111111" when X = 162 AND Y = 77 else
"111111111111" when X = 163 AND Y = 77 else
"111111111111" when X = 164 AND Y = 77 else
"111111111111" when X = 165 AND Y = 77 else
"111111111111" when X = 166 AND Y = 77 else
"111111111111" when X = 167 AND Y = 77 else
"111111111111" when X = 168 AND Y = 77 else
"111111111111" when X = 169 AND Y = 77 else
"111111111111" when X = 170 AND Y = 77 else
"111111111111" when X = 171 AND Y = 77 else
"111111111111" when X = 172 AND Y = 77 else
"111111111111" when X = 173 AND Y = 77 else
"111111111111" when X = 174 AND Y = 77 else
"111111111111" when X = 175 AND Y = 77 else
"111111111111" when X = 176 AND Y = 77 else
"111111111111" when X = 177 AND Y = 77 else
"111111111111" when X = 178 AND Y = 77 else
"111111111111" when X = 179 AND Y = 77 else
"111111111111" when X = 180 AND Y = 77 else
"111111111111" when X = 181 AND Y = 77 else
"111111111111" when X = 182 AND Y = 77 else
"111111111111" when X = 183 AND Y = 77 else
"111111111111" when X = 184 AND Y = 77 else
"111111111111" when X = 185 AND Y = 77 else
"111111111111" when X = 186 AND Y = 77 else
"111111111111" when X = 187 AND Y = 77 else
"111111111111" when X = 188 AND Y = 77 else
"111111111111" when X = 189 AND Y = 77 else
"111111111111" when X = 190 AND Y = 77 else
"111111111111" when X = 191 AND Y = 77 else
"111111111111" when X = 192 AND Y = 77 else
"111111111111" when X = 193 AND Y = 77 else
"111111111111" when X = 194 AND Y = 77 else
"111111111111" when X = 195 AND Y = 77 else
"111111111111" when X = 196 AND Y = 77 else
"111111111111" when X = 197 AND Y = 77 else
"111111111111" when X = 198 AND Y = 77 else
"111111111111" when X = 199 AND Y = 77 else
"111111111111" when X = 200 AND Y = 77 else
"111111111111" when X = 201 AND Y = 77 else
"111111111111" when X = 202 AND Y = 77 else
"111111111111" when X = 203 AND Y = 77 else
"111111111111" when X = 204 AND Y = 77 else
"111111111111" when X = 205 AND Y = 77 else
"111111111111" when X = 206 AND Y = 77 else
"111111111111" when X = 207 AND Y = 77 else
"111111111111" when X = 208 AND Y = 77 else
"111111111111" when X = 209 AND Y = 77 else
"111111111111" when X = 210 AND Y = 77 else
"111111111111" when X = 211 AND Y = 77 else
"111111111111" when X = 212 AND Y = 77 else
"111111111111" when X = 213 AND Y = 77 else
"111111111111" when X = 214 AND Y = 77 else
"111111111111" when X = 215 AND Y = 77 else
"111111111111" when X = 216 AND Y = 77 else
"111111111111" when X = 217 AND Y = 77 else
"111111111111" when X = 218 AND Y = 77 else
"111111111111" when X = 219 AND Y = 77 else
"111111111111" when X = 220 AND Y = 77 else
"111111111111" when X = 221 AND Y = 77 else
"111111111111" when X = 222 AND Y = 77 else
"111111111111" when X = 223 AND Y = 77 else
"111111111111" when X = 224 AND Y = 77 else
"111111111111" when X = 225 AND Y = 77 else
"111111111111" when X = 226 AND Y = 77 else
"111111111111" when X = 227 AND Y = 77 else
"111111111111" when X = 228 AND Y = 77 else
"111111111111" when X = 229 AND Y = 77 else
"111111111111" when X = 230 AND Y = 77 else
"111111111111" when X = 231 AND Y = 77 else
"111111111111" when X = 232 AND Y = 77 else
"111111111111" when X = 233 AND Y = 77 else
"111111111111" when X = 234 AND Y = 77 else
"111111111111" when X = 235 AND Y = 77 else
"111111111111" when X = 236 AND Y = 77 else
"111111111111" when X = 237 AND Y = 77 else
"111111111111" when X = 238 AND Y = 77 else
"111111111111" when X = 239 AND Y = 77 else
"111111111111" when X = 240 AND Y = 77 else
"111111111111" when X = 241 AND Y = 77 else
"111111111111" when X = 242 AND Y = 77 else
"111111111111" when X = 243 AND Y = 77 else
"111111111111" when X = 244 AND Y = 77 else
"111111111111" when X = 245 AND Y = 77 else
"111111111111" when X = 246 AND Y = 77 else
"111111111111" when X = 247 AND Y = 77 else
"111111111111" when X = 248 AND Y = 77 else
"111111111111" when X = 249 AND Y = 77 else
"111111111111" when X = 250 AND Y = 77 else
"111111111111" when X = 251 AND Y = 77 else
"111111111111" when X = 252 AND Y = 77 else
"111111111111" when X = 253 AND Y = 77 else
"111111111111" when X = 254 AND Y = 77 else
"111111111111" when X = 255 AND Y = 77 else
"111111111111" when X = 256 AND Y = 77 else
"111111111111" when X = 257 AND Y = 77 else
"111111111111" when X = 258 AND Y = 77 else
"111111111111" when X = 259 AND Y = 77 else
"111111111111" when X = 260 AND Y = 77 else
"111111111111" when X = 261 AND Y = 77 else
"111111111111" when X = 262 AND Y = 77 else
"111111111111" when X = 263 AND Y = 77 else
"111111111111" when X = 264 AND Y = 77 else
"110111011111" when X = 265 AND Y = 77 else
"110111011111" when X = 266 AND Y = 77 else
"110111011111" when X = 267 AND Y = 77 else
"110111011111" when X = 268 AND Y = 77 else
"110111011111" when X = 269 AND Y = 77 else
"110111011111" when X = 270 AND Y = 77 else
"110111011111" when X = 271 AND Y = 77 else
"110111011111" when X = 272 AND Y = 77 else
"110111011111" when X = 273 AND Y = 77 else
"110111011111" when X = 274 AND Y = 77 else
"110111011111" when X = 275 AND Y = 77 else
"110111011111" when X = 276 AND Y = 77 else
"110111011111" when X = 277 AND Y = 77 else
"110111011111" when X = 278 AND Y = 77 else
"110111011111" when X = 279 AND Y = 77 else
"000000000000" when X = 280 AND Y = 77 else
"000000000000" when X = 281 AND Y = 77 else
"000000000000" when X = 282 AND Y = 77 else
"000000000000" when X = 283 AND Y = 77 else
"000000000000" when X = 284 AND Y = 77 else
"000000000000" when X = 285 AND Y = 77 else
"000000000000" when X = 286 AND Y = 77 else
"000000000000" when X = 287 AND Y = 77 else
"000000000000" when X = 288 AND Y = 77 else
"000000000000" when X = 289 AND Y = 77 else
"000000000000" when X = 290 AND Y = 77 else
"000000000000" when X = 291 AND Y = 77 else
"000000000000" when X = 292 AND Y = 77 else
"000000000000" when X = 293 AND Y = 77 else
"000000000000" when X = 294 AND Y = 77 else
"000000000000" when X = 295 AND Y = 77 else
"000000000000" when X = 296 AND Y = 77 else
"000000000000" when X = 297 AND Y = 77 else
"000000000000" when X = 298 AND Y = 77 else
"000000000000" when X = 299 AND Y = 77 else
"000000000000" when X = 300 AND Y = 77 else
"000000000000" when X = 301 AND Y = 77 else
"000000000000" when X = 302 AND Y = 77 else
"000000000000" when X = 303 AND Y = 77 else
"000000000000" when X = 304 AND Y = 77 else
"000000000000" when X = 305 AND Y = 77 else
"000000000000" when X = 306 AND Y = 77 else
"000000000000" when X = 307 AND Y = 77 else
"000000000000" when X = 308 AND Y = 77 else
"000000000000" when X = 309 AND Y = 77 else
"000000000000" when X = 310 AND Y = 77 else
"000000000000" when X = 311 AND Y = 77 else
"000000000000" when X = 312 AND Y = 77 else
"000000000000" when X = 313 AND Y = 77 else
"000000000000" when X = 314 AND Y = 77 else
"000000000000" when X = 315 AND Y = 77 else
"000000000000" when X = 316 AND Y = 77 else
"000000000000" when X = 317 AND Y = 77 else
"000000000000" when X = 318 AND Y = 77 else
"000000000000" when X = 319 AND Y = 77 else
"000000000000" when X = 320 AND Y = 77 else
"000000000000" when X = 321 AND Y = 77 else
"000000000000" when X = 322 AND Y = 77 else
"000000000000" when X = 323 AND Y = 77 else
"000000000000" when X = 324 AND Y = 77 else
"100010011101" when X = 0 AND Y = 78 else
"100010011101" when X = 1 AND Y = 78 else
"100010011101" when X = 2 AND Y = 78 else
"100010011101" when X = 3 AND Y = 78 else
"100010011101" when X = 4 AND Y = 78 else
"100010011101" when X = 5 AND Y = 78 else
"100010011101" when X = 6 AND Y = 78 else
"100010011101" when X = 7 AND Y = 78 else
"100010011101" when X = 8 AND Y = 78 else
"100010011101" when X = 9 AND Y = 78 else
"100010011101" when X = 10 AND Y = 78 else
"100010011101" when X = 11 AND Y = 78 else
"100010011101" when X = 12 AND Y = 78 else
"100010011101" when X = 13 AND Y = 78 else
"100010011101" when X = 14 AND Y = 78 else
"100010011101" when X = 15 AND Y = 78 else
"100010011101" when X = 16 AND Y = 78 else
"100010011101" when X = 17 AND Y = 78 else
"100010011101" when X = 18 AND Y = 78 else
"100010011101" when X = 19 AND Y = 78 else
"100010011101" when X = 20 AND Y = 78 else
"100010011101" when X = 21 AND Y = 78 else
"100010011101" when X = 22 AND Y = 78 else
"100010011101" when X = 23 AND Y = 78 else
"100010011101" when X = 24 AND Y = 78 else
"100010011101" when X = 25 AND Y = 78 else
"100010011101" when X = 26 AND Y = 78 else
"100010011101" when X = 27 AND Y = 78 else
"100010011101" when X = 28 AND Y = 78 else
"100010011101" when X = 29 AND Y = 78 else
"110111011111" when X = 30 AND Y = 78 else
"110111011111" when X = 31 AND Y = 78 else
"110111011111" when X = 32 AND Y = 78 else
"110111011111" when X = 33 AND Y = 78 else
"110111011111" when X = 34 AND Y = 78 else
"110111011111" when X = 35 AND Y = 78 else
"110111011111" when X = 36 AND Y = 78 else
"110111011111" when X = 37 AND Y = 78 else
"110111011111" when X = 38 AND Y = 78 else
"110111011111" when X = 39 AND Y = 78 else
"110111011111" when X = 40 AND Y = 78 else
"110111011111" when X = 41 AND Y = 78 else
"110111011111" when X = 42 AND Y = 78 else
"110111011111" when X = 43 AND Y = 78 else
"110111011111" when X = 44 AND Y = 78 else
"110111011111" when X = 45 AND Y = 78 else
"110111011111" when X = 46 AND Y = 78 else
"110111011111" when X = 47 AND Y = 78 else
"110111011111" when X = 48 AND Y = 78 else
"110111011111" when X = 49 AND Y = 78 else
"110111011111" when X = 50 AND Y = 78 else
"110111011111" when X = 51 AND Y = 78 else
"110111011111" when X = 52 AND Y = 78 else
"110111011111" when X = 53 AND Y = 78 else
"110111011111" when X = 54 AND Y = 78 else
"110111011111" when X = 55 AND Y = 78 else
"110111011111" when X = 56 AND Y = 78 else
"110111011111" when X = 57 AND Y = 78 else
"110111011111" when X = 58 AND Y = 78 else
"110111011111" when X = 59 AND Y = 78 else
"110111011111" when X = 60 AND Y = 78 else
"110111011111" when X = 61 AND Y = 78 else
"110111011111" when X = 62 AND Y = 78 else
"110111011111" when X = 63 AND Y = 78 else
"110111011111" when X = 64 AND Y = 78 else
"110111011111" when X = 65 AND Y = 78 else
"110111011111" when X = 66 AND Y = 78 else
"110111011111" when X = 67 AND Y = 78 else
"110111011111" when X = 68 AND Y = 78 else
"110111011111" when X = 69 AND Y = 78 else
"110111011111" when X = 70 AND Y = 78 else
"110111011111" when X = 71 AND Y = 78 else
"110111011111" when X = 72 AND Y = 78 else
"110111011111" when X = 73 AND Y = 78 else
"110111011111" when X = 74 AND Y = 78 else
"110111011111" when X = 75 AND Y = 78 else
"110111011111" when X = 76 AND Y = 78 else
"110111011111" when X = 77 AND Y = 78 else
"110111011111" when X = 78 AND Y = 78 else
"110111011111" when X = 79 AND Y = 78 else
"110111011111" when X = 80 AND Y = 78 else
"110111011111" when X = 81 AND Y = 78 else
"110111011111" when X = 82 AND Y = 78 else
"110111011111" when X = 83 AND Y = 78 else
"110111011111" when X = 84 AND Y = 78 else
"110111011111" when X = 85 AND Y = 78 else
"110111011111" when X = 86 AND Y = 78 else
"110111011111" when X = 87 AND Y = 78 else
"110111011111" when X = 88 AND Y = 78 else
"110111011111" when X = 89 AND Y = 78 else
"110111011111" when X = 90 AND Y = 78 else
"110111011111" when X = 91 AND Y = 78 else
"110111011111" when X = 92 AND Y = 78 else
"110111011111" when X = 93 AND Y = 78 else
"110111011111" when X = 94 AND Y = 78 else
"110111011111" when X = 95 AND Y = 78 else
"110111011111" when X = 96 AND Y = 78 else
"110111011111" when X = 97 AND Y = 78 else
"110111011111" when X = 98 AND Y = 78 else
"110111011111" when X = 99 AND Y = 78 else
"110111011111" when X = 100 AND Y = 78 else
"110111011111" when X = 101 AND Y = 78 else
"110111011111" when X = 102 AND Y = 78 else
"110111011111" when X = 103 AND Y = 78 else
"110111011111" when X = 104 AND Y = 78 else
"110111011111" when X = 105 AND Y = 78 else
"110111011111" when X = 106 AND Y = 78 else
"110111011111" when X = 107 AND Y = 78 else
"110111011111" when X = 108 AND Y = 78 else
"110111011111" when X = 109 AND Y = 78 else
"111111111111" when X = 110 AND Y = 78 else
"111111111111" when X = 111 AND Y = 78 else
"111111111111" when X = 112 AND Y = 78 else
"111111111111" when X = 113 AND Y = 78 else
"111111111111" when X = 114 AND Y = 78 else
"111111111111" when X = 115 AND Y = 78 else
"111111111111" when X = 116 AND Y = 78 else
"111111111111" when X = 117 AND Y = 78 else
"111111111111" when X = 118 AND Y = 78 else
"111111111111" when X = 119 AND Y = 78 else
"111111111111" when X = 120 AND Y = 78 else
"111111111111" when X = 121 AND Y = 78 else
"111111111111" when X = 122 AND Y = 78 else
"111111111111" when X = 123 AND Y = 78 else
"111111111111" when X = 124 AND Y = 78 else
"111111111111" when X = 125 AND Y = 78 else
"111111111111" when X = 126 AND Y = 78 else
"111111111111" when X = 127 AND Y = 78 else
"111111111111" when X = 128 AND Y = 78 else
"111111111111" when X = 129 AND Y = 78 else
"111111111111" when X = 130 AND Y = 78 else
"111111111111" when X = 131 AND Y = 78 else
"111111111111" when X = 132 AND Y = 78 else
"111111111111" when X = 133 AND Y = 78 else
"111111111111" when X = 134 AND Y = 78 else
"111111111111" when X = 135 AND Y = 78 else
"111111111111" when X = 136 AND Y = 78 else
"111111111111" when X = 137 AND Y = 78 else
"111111111111" when X = 138 AND Y = 78 else
"111111111111" when X = 139 AND Y = 78 else
"111111111111" when X = 140 AND Y = 78 else
"111111111111" when X = 141 AND Y = 78 else
"111111111111" when X = 142 AND Y = 78 else
"111111111111" when X = 143 AND Y = 78 else
"111111111111" when X = 144 AND Y = 78 else
"111111111111" when X = 145 AND Y = 78 else
"111111111111" when X = 146 AND Y = 78 else
"111111111111" when X = 147 AND Y = 78 else
"111111111111" when X = 148 AND Y = 78 else
"111111111111" when X = 149 AND Y = 78 else
"111111111111" when X = 150 AND Y = 78 else
"111111111111" when X = 151 AND Y = 78 else
"111111111111" when X = 152 AND Y = 78 else
"111111111111" when X = 153 AND Y = 78 else
"111111111111" when X = 154 AND Y = 78 else
"111111111111" when X = 155 AND Y = 78 else
"111111111111" when X = 156 AND Y = 78 else
"111111111111" when X = 157 AND Y = 78 else
"111111111111" when X = 158 AND Y = 78 else
"111111111111" when X = 159 AND Y = 78 else
"111111111111" when X = 160 AND Y = 78 else
"111111111111" when X = 161 AND Y = 78 else
"111111111111" when X = 162 AND Y = 78 else
"111111111111" when X = 163 AND Y = 78 else
"111111111111" when X = 164 AND Y = 78 else
"111111111111" when X = 165 AND Y = 78 else
"111111111111" when X = 166 AND Y = 78 else
"111111111111" when X = 167 AND Y = 78 else
"111111111111" when X = 168 AND Y = 78 else
"111111111111" when X = 169 AND Y = 78 else
"111111111111" when X = 170 AND Y = 78 else
"111111111111" when X = 171 AND Y = 78 else
"111111111111" when X = 172 AND Y = 78 else
"111111111111" when X = 173 AND Y = 78 else
"111111111111" when X = 174 AND Y = 78 else
"111111111111" when X = 175 AND Y = 78 else
"111111111111" when X = 176 AND Y = 78 else
"111111111111" when X = 177 AND Y = 78 else
"111111111111" when X = 178 AND Y = 78 else
"111111111111" when X = 179 AND Y = 78 else
"111111111111" when X = 180 AND Y = 78 else
"111111111111" when X = 181 AND Y = 78 else
"111111111111" when X = 182 AND Y = 78 else
"111111111111" when X = 183 AND Y = 78 else
"111111111111" when X = 184 AND Y = 78 else
"111111111111" when X = 185 AND Y = 78 else
"111111111111" when X = 186 AND Y = 78 else
"111111111111" when X = 187 AND Y = 78 else
"111111111111" when X = 188 AND Y = 78 else
"111111111111" when X = 189 AND Y = 78 else
"111111111111" when X = 190 AND Y = 78 else
"111111111111" when X = 191 AND Y = 78 else
"111111111111" when X = 192 AND Y = 78 else
"111111111111" when X = 193 AND Y = 78 else
"111111111111" when X = 194 AND Y = 78 else
"111111111111" when X = 195 AND Y = 78 else
"111111111111" when X = 196 AND Y = 78 else
"111111111111" when X = 197 AND Y = 78 else
"111111111111" when X = 198 AND Y = 78 else
"111111111111" when X = 199 AND Y = 78 else
"111111111111" when X = 200 AND Y = 78 else
"111111111111" when X = 201 AND Y = 78 else
"111111111111" when X = 202 AND Y = 78 else
"111111111111" when X = 203 AND Y = 78 else
"111111111111" when X = 204 AND Y = 78 else
"111111111111" when X = 205 AND Y = 78 else
"111111111111" when X = 206 AND Y = 78 else
"111111111111" when X = 207 AND Y = 78 else
"111111111111" when X = 208 AND Y = 78 else
"111111111111" when X = 209 AND Y = 78 else
"111111111111" when X = 210 AND Y = 78 else
"111111111111" when X = 211 AND Y = 78 else
"111111111111" when X = 212 AND Y = 78 else
"111111111111" when X = 213 AND Y = 78 else
"111111111111" when X = 214 AND Y = 78 else
"111111111111" when X = 215 AND Y = 78 else
"111111111111" when X = 216 AND Y = 78 else
"111111111111" when X = 217 AND Y = 78 else
"111111111111" when X = 218 AND Y = 78 else
"111111111111" when X = 219 AND Y = 78 else
"111111111111" when X = 220 AND Y = 78 else
"111111111111" when X = 221 AND Y = 78 else
"111111111111" when X = 222 AND Y = 78 else
"111111111111" when X = 223 AND Y = 78 else
"111111111111" when X = 224 AND Y = 78 else
"111111111111" when X = 225 AND Y = 78 else
"111111111111" when X = 226 AND Y = 78 else
"111111111111" when X = 227 AND Y = 78 else
"111111111111" when X = 228 AND Y = 78 else
"111111111111" when X = 229 AND Y = 78 else
"111111111111" when X = 230 AND Y = 78 else
"111111111111" when X = 231 AND Y = 78 else
"111111111111" when X = 232 AND Y = 78 else
"111111111111" when X = 233 AND Y = 78 else
"111111111111" when X = 234 AND Y = 78 else
"111111111111" when X = 235 AND Y = 78 else
"111111111111" when X = 236 AND Y = 78 else
"111111111111" when X = 237 AND Y = 78 else
"111111111111" when X = 238 AND Y = 78 else
"111111111111" when X = 239 AND Y = 78 else
"111111111111" when X = 240 AND Y = 78 else
"111111111111" when X = 241 AND Y = 78 else
"111111111111" when X = 242 AND Y = 78 else
"111111111111" when X = 243 AND Y = 78 else
"111111111111" when X = 244 AND Y = 78 else
"111111111111" when X = 245 AND Y = 78 else
"111111111111" when X = 246 AND Y = 78 else
"111111111111" when X = 247 AND Y = 78 else
"111111111111" when X = 248 AND Y = 78 else
"111111111111" when X = 249 AND Y = 78 else
"111111111111" when X = 250 AND Y = 78 else
"111111111111" when X = 251 AND Y = 78 else
"111111111111" when X = 252 AND Y = 78 else
"111111111111" when X = 253 AND Y = 78 else
"111111111111" when X = 254 AND Y = 78 else
"111111111111" when X = 255 AND Y = 78 else
"111111111111" when X = 256 AND Y = 78 else
"111111111111" when X = 257 AND Y = 78 else
"111111111111" when X = 258 AND Y = 78 else
"111111111111" when X = 259 AND Y = 78 else
"111111111111" when X = 260 AND Y = 78 else
"111111111111" when X = 261 AND Y = 78 else
"111111111111" when X = 262 AND Y = 78 else
"111111111111" when X = 263 AND Y = 78 else
"111111111111" when X = 264 AND Y = 78 else
"110111011111" when X = 265 AND Y = 78 else
"110111011111" when X = 266 AND Y = 78 else
"110111011111" when X = 267 AND Y = 78 else
"110111011111" when X = 268 AND Y = 78 else
"110111011111" when X = 269 AND Y = 78 else
"110111011111" when X = 270 AND Y = 78 else
"110111011111" when X = 271 AND Y = 78 else
"110111011111" when X = 272 AND Y = 78 else
"110111011111" when X = 273 AND Y = 78 else
"110111011111" when X = 274 AND Y = 78 else
"110111011111" when X = 275 AND Y = 78 else
"110111011111" when X = 276 AND Y = 78 else
"110111011111" when X = 277 AND Y = 78 else
"110111011111" when X = 278 AND Y = 78 else
"110111011111" when X = 279 AND Y = 78 else
"000000000000" when X = 280 AND Y = 78 else
"000000000000" when X = 281 AND Y = 78 else
"000000000000" when X = 282 AND Y = 78 else
"000000000000" when X = 283 AND Y = 78 else
"000000000000" when X = 284 AND Y = 78 else
"000000000000" when X = 285 AND Y = 78 else
"000000000000" when X = 286 AND Y = 78 else
"000000000000" when X = 287 AND Y = 78 else
"000000000000" when X = 288 AND Y = 78 else
"000000000000" when X = 289 AND Y = 78 else
"000000000000" when X = 290 AND Y = 78 else
"000000000000" when X = 291 AND Y = 78 else
"000000000000" when X = 292 AND Y = 78 else
"000000000000" when X = 293 AND Y = 78 else
"000000000000" when X = 294 AND Y = 78 else
"000000000000" when X = 295 AND Y = 78 else
"000000000000" when X = 296 AND Y = 78 else
"000000000000" when X = 297 AND Y = 78 else
"000000000000" when X = 298 AND Y = 78 else
"000000000000" when X = 299 AND Y = 78 else
"000000000000" when X = 300 AND Y = 78 else
"000000000000" when X = 301 AND Y = 78 else
"000000000000" when X = 302 AND Y = 78 else
"000000000000" when X = 303 AND Y = 78 else
"000000000000" when X = 304 AND Y = 78 else
"000000000000" when X = 305 AND Y = 78 else
"000000000000" when X = 306 AND Y = 78 else
"000000000000" when X = 307 AND Y = 78 else
"000000000000" when X = 308 AND Y = 78 else
"000000000000" when X = 309 AND Y = 78 else
"000000000000" when X = 310 AND Y = 78 else
"000000000000" when X = 311 AND Y = 78 else
"000000000000" when X = 312 AND Y = 78 else
"000000000000" when X = 313 AND Y = 78 else
"000000000000" when X = 314 AND Y = 78 else
"000000000000" when X = 315 AND Y = 78 else
"000000000000" when X = 316 AND Y = 78 else
"000000000000" when X = 317 AND Y = 78 else
"000000000000" when X = 318 AND Y = 78 else
"000000000000" when X = 319 AND Y = 78 else
"000000000000" when X = 320 AND Y = 78 else
"000000000000" when X = 321 AND Y = 78 else
"000000000000" when X = 322 AND Y = 78 else
"000000000000" when X = 323 AND Y = 78 else
"000000000000" when X = 324 AND Y = 78 else
"100010011101" when X = 0 AND Y = 79 else
"100010011101" when X = 1 AND Y = 79 else
"100010011101" when X = 2 AND Y = 79 else
"100010011101" when X = 3 AND Y = 79 else
"100010011101" when X = 4 AND Y = 79 else
"100010011101" when X = 5 AND Y = 79 else
"100010011101" when X = 6 AND Y = 79 else
"100010011101" when X = 7 AND Y = 79 else
"100010011101" when X = 8 AND Y = 79 else
"100010011101" when X = 9 AND Y = 79 else
"100010011101" when X = 10 AND Y = 79 else
"100010011101" when X = 11 AND Y = 79 else
"100010011101" when X = 12 AND Y = 79 else
"100010011101" when X = 13 AND Y = 79 else
"100010011101" when X = 14 AND Y = 79 else
"100010011101" when X = 15 AND Y = 79 else
"100010011101" when X = 16 AND Y = 79 else
"100010011101" when X = 17 AND Y = 79 else
"100010011101" when X = 18 AND Y = 79 else
"100010011101" when X = 19 AND Y = 79 else
"100010011101" when X = 20 AND Y = 79 else
"100010011101" when X = 21 AND Y = 79 else
"100010011101" when X = 22 AND Y = 79 else
"100010011101" when X = 23 AND Y = 79 else
"100010011101" when X = 24 AND Y = 79 else
"100010011101" when X = 25 AND Y = 79 else
"100010011101" when X = 26 AND Y = 79 else
"100010011101" when X = 27 AND Y = 79 else
"100010011101" when X = 28 AND Y = 79 else
"100010011101" when X = 29 AND Y = 79 else
"110111011111" when X = 30 AND Y = 79 else
"110111011111" when X = 31 AND Y = 79 else
"110111011111" when X = 32 AND Y = 79 else
"110111011111" when X = 33 AND Y = 79 else
"110111011111" when X = 34 AND Y = 79 else
"110111011111" when X = 35 AND Y = 79 else
"110111011111" when X = 36 AND Y = 79 else
"110111011111" when X = 37 AND Y = 79 else
"110111011111" when X = 38 AND Y = 79 else
"110111011111" when X = 39 AND Y = 79 else
"110111011111" when X = 40 AND Y = 79 else
"110111011111" when X = 41 AND Y = 79 else
"110111011111" when X = 42 AND Y = 79 else
"110111011111" when X = 43 AND Y = 79 else
"110111011111" when X = 44 AND Y = 79 else
"110111011111" when X = 45 AND Y = 79 else
"110111011111" when X = 46 AND Y = 79 else
"110111011111" when X = 47 AND Y = 79 else
"110111011111" when X = 48 AND Y = 79 else
"110111011111" when X = 49 AND Y = 79 else
"110111011111" when X = 50 AND Y = 79 else
"110111011111" when X = 51 AND Y = 79 else
"110111011111" when X = 52 AND Y = 79 else
"110111011111" when X = 53 AND Y = 79 else
"110111011111" when X = 54 AND Y = 79 else
"110111011111" when X = 55 AND Y = 79 else
"110111011111" when X = 56 AND Y = 79 else
"110111011111" when X = 57 AND Y = 79 else
"110111011111" when X = 58 AND Y = 79 else
"110111011111" when X = 59 AND Y = 79 else
"110111011111" when X = 60 AND Y = 79 else
"110111011111" when X = 61 AND Y = 79 else
"110111011111" when X = 62 AND Y = 79 else
"110111011111" when X = 63 AND Y = 79 else
"110111011111" when X = 64 AND Y = 79 else
"110111011111" when X = 65 AND Y = 79 else
"110111011111" when X = 66 AND Y = 79 else
"110111011111" when X = 67 AND Y = 79 else
"110111011111" when X = 68 AND Y = 79 else
"110111011111" when X = 69 AND Y = 79 else
"110111011111" when X = 70 AND Y = 79 else
"110111011111" when X = 71 AND Y = 79 else
"110111011111" when X = 72 AND Y = 79 else
"110111011111" when X = 73 AND Y = 79 else
"110111011111" when X = 74 AND Y = 79 else
"110111011111" when X = 75 AND Y = 79 else
"110111011111" when X = 76 AND Y = 79 else
"110111011111" when X = 77 AND Y = 79 else
"110111011111" when X = 78 AND Y = 79 else
"110111011111" when X = 79 AND Y = 79 else
"110111011111" when X = 80 AND Y = 79 else
"110111011111" when X = 81 AND Y = 79 else
"110111011111" when X = 82 AND Y = 79 else
"110111011111" when X = 83 AND Y = 79 else
"110111011111" when X = 84 AND Y = 79 else
"110111011111" when X = 85 AND Y = 79 else
"110111011111" when X = 86 AND Y = 79 else
"110111011111" when X = 87 AND Y = 79 else
"110111011111" when X = 88 AND Y = 79 else
"110111011111" when X = 89 AND Y = 79 else
"110111011111" when X = 90 AND Y = 79 else
"110111011111" when X = 91 AND Y = 79 else
"110111011111" when X = 92 AND Y = 79 else
"110111011111" when X = 93 AND Y = 79 else
"110111011111" when X = 94 AND Y = 79 else
"110111011111" when X = 95 AND Y = 79 else
"110111011111" when X = 96 AND Y = 79 else
"110111011111" when X = 97 AND Y = 79 else
"110111011111" when X = 98 AND Y = 79 else
"110111011111" when X = 99 AND Y = 79 else
"110111011111" when X = 100 AND Y = 79 else
"110111011111" when X = 101 AND Y = 79 else
"110111011111" when X = 102 AND Y = 79 else
"110111011111" when X = 103 AND Y = 79 else
"110111011111" when X = 104 AND Y = 79 else
"110111011111" when X = 105 AND Y = 79 else
"110111011111" when X = 106 AND Y = 79 else
"110111011111" when X = 107 AND Y = 79 else
"110111011111" when X = 108 AND Y = 79 else
"110111011111" when X = 109 AND Y = 79 else
"111111111111" when X = 110 AND Y = 79 else
"111111111111" when X = 111 AND Y = 79 else
"111111111111" when X = 112 AND Y = 79 else
"111111111111" when X = 113 AND Y = 79 else
"111111111111" when X = 114 AND Y = 79 else
"111111111111" when X = 115 AND Y = 79 else
"111111111111" when X = 116 AND Y = 79 else
"111111111111" when X = 117 AND Y = 79 else
"111111111111" when X = 118 AND Y = 79 else
"111111111111" when X = 119 AND Y = 79 else
"111111111111" when X = 120 AND Y = 79 else
"111111111111" when X = 121 AND Y = 79 else
"111111111111" when X = 122 AND Y = 79 else
"111111111111" when X = 123 AND Y = 79 else
"111111111111" when X = 124 AND Y = 79 else
"111111111111" when X = 125 AND Y = 79 else
"111111111111" when X = 126 AND Y = 79 else
"111111111111" when X = 127 AND Y = 79 else
"111111111111" when X = 128 AND Y = 79 else
"111111111111" when X = 129 AND Y = 79 else
"111111111111" when X = 130 AND Y = 79 else
"111111111111" when X = 131 AND Y = 79 else
"111111111111" when X = 132 AND Y = 79 else
"111111111111" when X = 133 AND Y = 79 else
"111111111111" when X = 134 AND Y = 79 else
"111111111111" when X = 135 AND Y = 79 else
"111111111111" when X = 136 AND Y = 79 else
"111111111111" when X = 137 AND Y = 79 else
"111111111111" when X = 138 AND Y = 79 else
"111111111111" when X = 139 AND Y = 79 else
"111111111111" when X = 140 AND Y = 79 else
"111111111111" when X = 141 AND Y = 79 else
"111111111111" when X = 142 AND Y = 79 else
"111111111111" when X = 143 AND Y = 79 else
"111111111111" when X = 144 AND Y = 79 else
"111111111111" when X = 145 AND Y = 79 else
"111111111111" when X = 146 AND Y = 79 else
"111111111111" when X = 147 AND Y = 79 else
"111111111111" when X = 148 AND Y = 79 else
"111111111111" when X = 149 AND Y = 79 else
"111111111111" when X = 150 AND Y = 79 else
"111111111111" when X = 151 AND Y = 79 else
"111111111111" when X = 152 AND Y = 79 else
"111111111111" when X = 153 AND Y = 79 else
"111111111111" when X = 154 AND Y = 79 else
"111111111111" when X = 155 AND Y = 79 else
"111111111111" when X = 156 AND Y = 79 else
"111111111111" when X = 157 AND Y = 79 else
"111111111111" when X = 158 AND Y = 79 else
"111111111111" when X = 159 AND Y = 79 else
"111111111111" when X = 160 AND Y = 79 else
"111111111111" when X = 161 AND Y = 79 else
"111111111111" when X = 162 AND Y = 79 else
"111111111111" when X = 163 AND Y = 79 else
"111111111111" when X = 164 AND Y = 79 else
"111111111111" when X = 165 AND Y = 79 else
"111111111111" when X = 166 AND Y = 79 else
"111111111111" when X = 167 AND Y = 79 else
"111111111111" when X = 168 AND Y = 79 else
"111111111111" when X = 169 AND Y = 79 else
"111111111111" when X = 170 AND Y = 79 else
"111111111111" when X = 171 AND Y = 79 else
"111111111111" when X = 172 AND Y = 79 else
"111111111111" when X = 173 AND Y = 79 else
"111111111111" when X = 174 AND Y = 79 else
"111111111111" when X = 175 AND Y = 79 else
"111111111111" when X = 176 AND Y = 79 else
"111111111111" when X = 177 AND Y = 79 else
"111111111111" when X = 178 AND Y = 79 else
"111111111111" when X = 179 AND Y = 79 else
"111111111111" when X = 180 AND Y = 79 else
"111111111111" when X = 181 AND Y = 79 else
"111111111111" when X = 182 AND Y = 79 else
"111111111111" when X = 183 AND Y = 79 else
"111111111111" when X = 184 AND Y = 79 else
"111111111111" when X = 185 AND Y = 79 else
"111111111111" when X = 186 AND Y = 79 else
"111111111111" when X = 187 AND Y = 79 else
"111111111111" when X = 188 AND Y = 79 else
"111111111111" when X = 189 AND Y = 79 else
"111111111111" when X = 190 AND Y = 79 else
"111111111111" when X = 191 AND Y = 79 else
"111111111111" when X = 192 AND Y = 79 else
"111111111111" when X = 193 AND Y = 79 else
"111111111111" when X = 194 AND Y = 79 else
"111111111111" when X = 195 AND Y = 79 else
"111111111111" when X = 196 AND Y = 79 else
"111111111111" when X = 197 AND Y = 79 else
"111111111111" when X = 198 AND Y = 79 else
"111111111111" when X = 199 AND Y = 79 else
"111111111111" when X = 200 AND Y = 79 else
"111111111111" when X = 201 AND Y = 79 else
"111111111111" when X = 202 AND Y = 79 else
"111111111111" when X = 203 AND Y = 79 else
"111111111111" when X = 204 AND Y = 79 else
"111111111111" when X = 205 AND Y = 79 else
"111111111111" when X = 206 AND Y = 79 else
"111111111111" when X = 207 AND Y = 79 else
"111111111111" when X = 208 AND Y = 79 else
"111111111111" when X = 209 AND Y = 79 else
"111111111111" when X = 210 AND Y = 79 else
"111111111111" when X = 211 AND Y = 79 else
"111111111111" when X = 212 AND Y = 79 else
"111111111111" when X = 213 AND Y = 79 else
"111111111111" when X = 214 AND Y = 79 else
"111111111111" when X = 215 AND Y = 79 else
"111111111111" when X = 216 AND Y = 79 else
"111111111111" when X = 217 AND Y = 79 else
"111111111111" when X = 218 AND Y = 79 else
"111111111111" when X = 219 AND Y = 79 else
"111111111111" when X = 220 AND Y = 79 else
"111111111111" when X = 221 AND Y = 79 else
"111111111111" when X = 222 AND Y = 79 else
"111111111111" when X = 223 AND Y = 79 else
"111111111111" when X = 224 AND Y = 79 else
"111111111111" when X = 225 AND Y = 79 else
"111111111111" when X = 226 AND Y = 79 else
"111111111111" when X = 227 AND Y = 79 else
"111111111111" when X = 228 AND Y = 79 else
"111111111111" when X = 229 AND Y = 79 else
"111111111111" when X = 230 AND Y = 79 else
"111111111111" when X = 231 AND Y = 79 else
"111111111111" when X = 232 AND Y = 79 else
"111111111111" when X = 233 AND Y = 79 else
"111111111111" when X = 234 AND Y = 79 else
"111111111111" when X = 235 AND Y = 79 else
"111111111111" when X = 236 AND Y = 79 else
"111111111111" when X = 237 AND Y = 79 else
"111111111111" when X = 238 AND Y = 79 else
"111111111111" when X = 239 AND Y = 79 else
"111111111111" when X = 240 AND Y = 79 else
"111111111111" when X = 241 AND Y = 79 else
"111111111111" when X = 242 AND Y = 79 else
"111111111111" when X = 243 AND Y = 79 else
"111111111111" when X = 244 AND Y = 79 else
"111111111111" when X = 245 AND Y = 79 else
"111111111111" when X = 246 AND Y = 79 else
"111111111111" when X = 247 AND Y = 79 else
"111111111111" when X = 248 AND Y = 79 else
"111111111111" when X = 249 AND Y = 79 else
"111111111111" when X = 250 AND Y = 79 else
"111111111111" when X = 251 AND Y = 79 else
"111111111111" when X = 252 AND Y = 79 else
"111111111111" when X = 253 AND Y = 79 else
"111111111111" when X = 254 AND Y = 79 else
"111111111111" when X = 255 AND Y = 79 else
"111111111111" when X = 256 AND Y = 79 else
"111111111111" when X = 257 AND Y = 79 else
"111111111111" when X = 258 AND Y = 79 else
"111111111111" when X = 259 AND Y = 79 else
"111111111111" when X = 260 AND Y = 79 else
"111111111111" when X = 261 AND Y = 79 else
"111111111111" when X = 262 AND Y = 79 else
"111111111111" when X = 263 AND Y = 79 else
"111111111111" when X = 264 AND Y = 79 else
"110111011111" when X = 265 AND Y = 79 else
"110111011111" when X = 266 AND Y = 79 else
"110111011111" when X = 267 AND Y = 79 else
"110111011111" when X = 268 AND Y = 79 else
"110111011111" when X = 269 AND Y = 79 else
"110111011111" when X = 270 AND Y = 79 else
"110111011111" when X = 271 AND Y = 79 else
"110111011111" when X = 272 AND Y = 79 else
"110111011111" when X = 273 AND Y = 79 else
"110111011111" when X = 274 AND Y = 79 else
"110111011111" when X = 275 AND Y = 79 else
"110111011111" when X = 276 AND Y = 79 else
"110111011111" when X = 277 AND Y = 79 else
"110111011111" when X = 278 AND Y = 79 else
"110111011111" when X = 279 AND Y = 79 else
"000000000000" when X = 280 AND Y = 79 else
"000000000000" when X = 281 AND Y = 79 else
"000000000000" when X = 282 AND Y = 79 else
"000000000000" when X = 283 AND Y = 79 else
"000000000000" when X = 284 AND Y = 79 else
"000000000000" when X = 285 AND Y = 79 else
"000000000000" when X = 286 AND Y = 79 else
"000000000000" when X = 287 AND Y = 79 else
"000000000000" when X = 288 AND Y = 79 else
"000000000000" when X = 289 AND Y = 79 else
"000000000000" when X = 290 AND Y = 79 else
"000000000000" when X = 291 AND Y = 79 else
"000000000000" when X = 292 AND Y = 79 else
"000000000000" when X = 293 AND Y = 79 else
"000000000000" when X = 294 AND Y = 79 else
"000000000000" when X = 295 AND Y = 79 else
"000000000000" when X = 296 AND Y = 79 else
"000000000000" when X = 297 AND Y = 79 else
"000000000000" when X = 298 AND Y = 79 else
"000000000000" when X = 299 AND Y = 79 else
"000000000000" when X = 300 AND Y = 79 else
"000000000000" when X = 301 AND Y = 79 else
"000000000000" when X = 302 AND Y = 79 else
"000000000000" when X = 303 AND Y = 79 else
"000000000000" when X = 304 AND Y = 79 else
"000000000000" when X = 305 AND Y = 79 else
"000000000000" when X = 306 AND Y = 79 else
"000000000000" when X = 307 AND Y = 79 else
"000000000000" when X = 308 AND Y = 79 else
"000000000000" when X = 309 AND Y = 79 else
"000000000000" when X = 310 AND Y = 79 else
"000000000000" when X = 311 AND Y = 79 else
"000000000000" when X = 312 AND Y = 79 else
"000000000000" when X = 313 AND Y = 79 else
"000000000000" when X = 314 AND Y = 79 else
"000000000000" when X = 315 AND Y = 79 else
"000000000000" when X = 316 AND Y = 79 else
"000000000000" when X = 317 AND Y = 79 else
"000000000000" when X = 318 AND Y = 79 else
"000000000000" when X = 319 AND Y = 79 else
"000000000000" when X = 320 AND Y = 79 else
"000000000000" when X = 321 AND Y = 79 else
"000000000000" when X = 322 AND Y = 79 else
"000000000000" when X = 323 AND Y = 79 else
"000000000000" when X = 324 AND Y = 79 else
"100010011101" when X = 0 AND Y = 80 else
"100010011101" when X = 1 AND Y = 80 else
"100010011101" when X = 2 AND Y = 80 else
"100010011101" when X = 3 AND Y = 80 else
"100010011101" when X = 4 AND Y = 80 else
"100010011101" when X = 5 AND Y = 80 else
"100010011101" when X = 6 AND Y = 80 else
"100010011101" when X = 7 AND Y = 80 else
"100010011101" when X = 8 AND Y = 80 else
"100010011101" when X = 9 AND Y = 80 else
"100010011101" when X = 10 AND Y = 80 else
"100010011101" when X = 11 AND Y = 80 else
"100010011101" when X = 12 AND Y = 80 else
"100010011101" when X = 13 AND Y = 80 else
"100010011101" when X = 14 AND Y = 80 else
"100010011101" when X = 15 AND Y = 80 else
"100010011101" when X = 16 AND Y = 80 else
"100010011101" when X = 17 AND Y = 80 else
"100010011101" when X = 18 AND Y = 80 else
"100010011101" when X = 19 AND Y = 80 else
"100010011101" when X = 20 AND Y = 80 else
"100010011101" when X = 21 AND Y = 80 else
"100010011101" when X = 22 AND Y = 80 else
"100010011101" when X = 23 AND Y = 80 else
"100010011101" when X = 24 AND Y = 80 else
"100010011101" when X = 25 AND Y = 80 else
"100010011101" when X = 26 AND Y = 80 else
"100010011101" when X = 27 AND Y = 80 else
"100010011101" when X = 28 AND Y = 80 else
"100010011101" when X = 29 AND Y = 80 else
"110111011111" when X = 30 AND Y = 80 else
"110111011111" when X = 31 AND Y = 80 else
"110111011111" when X = 32 AND Y = 80 else
"110111011111" when X = 33 AND Y = 80 else
"110111011111" when X = 34 AND Y = 80 else
"110111011111" when X = 35 AND Y = 80 else
"110111011111" when X = 36 AND Y = 80 else
"110111011111" when X = 37 AND Y = 80 else
"110111011111" when X = 38 AND Y = 80 else
"110111011111" when X = 39 AND Y = 80 else
"110111011111" when X = 40 AND Y = 80 else
"110111011111" when X = 41 AND Y = 80 else
"110111011111" when X = 42 AND Y = 80 else
"110111011111" when X = 43 AND Y = 80 else
"110111011111" when X = 44 AND Y = 80 else
"110111011111" when X = 45 AND Y = 80 else
"110111011111" when X = 46 AND Y = 80 else
"110111011111" when X = 47 AND Y = 80 else
"110111011111" when X = 48 AND Y = 80 else
"110111011111" when X = 49 AND Y = 80 else
"110111011111" when X = 50 AND Y = 80 else
"110111011111" when X = 51 AND Y = 80 else
"110111011111" when X = 52 AND Y = 80 else
"110111011111" when X = 53 AND Y = 80 else
"110111011111" when X = 54 AND Y = 80 else
"110111011111" when X = 55 AND Y = 80 else
"110111011111" when X = 56 AND Y = 80 else
"110111011111" when X = 57 AND Y = 80 else
"110111011111" when X = 58 AND Y = 80 else
"110111011111" when X = 59 AND Y = 80 else
"110111011111" when X = 60 AND Y = 80 else
"110111011111" when X = 61 AND Y = 80 else
"110111011111" when X = 62 AND Y = 80 else
"110111011111" when X = 63 AND Y = 80 else
"110111011111" when X = 64 AND Y = 80 else
"110111011111" when X = 65 AND Y = 80 else
"110111011111" when X = 66 AND Y = 80 else
"110111011111" when X = 67 AND Y = 80 else
"110111011111" when X = 68 AND Y = 80 else
"110111011111" when X = 69 AND Y = 80 else
"110111011111" when X = 70 AND Y = 80 else
"110111011111" when X = 71 AND Y = 80 else
"110111011111" when X = 72 AND Y = 80 else
"110111011111" when X = 73 AND Y = 80 else
"110111011111" when X = 74 AND Y = 80 else
"110111011111" when X = 75 AND Y = 80 else
"110111011111" when X = 76 AND Y = 80 else
"110111011111" when X = 77 AND Y = 80 else
"110111011111" when X = 78 AND Y = 80 else
"110111011111" when X = 79 AND Y = 80 else
"110111011111" when X = 80 AND Y = 80 else
"110111011111" when X = 81 AND Y = 80 else
"110111011111" when X = 82 AND Y = 80 else
"110111011111" when X = 83 AND Y = 80 else
"110111011111" when X = 84 AND Y = 80 else
"110111011111" when X = 85 AND Y = 80 else
"110111011111" when X = 86 AND Y = 80 else
"110111011111" when X = 87 AND Y = 80 else
"110111011111" when X = 88 AND Y = 80 else
"110111011111" when X = 89 AND Y = 80 else
"110111011111" when X = 90 AND Y = 80 else
"110111011111" when X = 91 AND Y = 80 else
"110111011111" when X = 92 AND Y = 80 else
"110111011111" when X = 93 AND Y = 80 else
"110111011111" when X = 94 AND Y = 80 else
"110111011111" when X = 95 AND Y = 80 else
"110111011111" when X = 96 AND Y = 80 else
"110111011111" when X = 97 AND Y = 80 else
"110111011111" when X = 98 AND Y = 80 else
"110111011111" when X = 99 AND Y = 80 else
"110111011111" when X = 100 AND Y = 80 else
"110111011111" when X = 101 AND Y = 80 else
"110111011111" when X = 102 AND Y = 80 else
"110111011111" when X = 103 AND Y = 80 else
"110111011111" when X = 104 AND Y = 80 else
"111111111111" when X = 105 AND Y = 80 else
"111111111111" when X = 106 AND Y = 80 else
"111111111111" when X = 107 AND Y = 80 else
"111111111111" when X = 108 AND Y = 80 else
"111111111111" when X = 109 AND Y = 80 else
"111111111111" when X = 110 AND Y = 80 else
"111111111111" when X = 111 AND Y = 80 else
"111111111111" when X = 112 AND Y = 80 else
"111111111111" when X = 113 AND Y = 80 else
"111111111111" when X = 114 AND Y = 80 else
"111111111111" when X = 115 AND Y = 80 else
"111111111111" when X = 116 AND Y = 80 else
"111111111111" when X = 117 AND Y = 80 else
"111111111111" when X = 118 AND Y = 80 else
"111111111111" when X = 119 AND Y = 80 else
"111111111111" when X = 120 AND Y = 80 else
"111111111111" when X = 121 AND Y = 80 else
"111111111111" when X = 122 AND Y = 80 else
"111111111111" when X = 123 AND Y = 80 else
"111111111111" when X = 124 AND Y = 80 else
"111111111111" when X = 125 AND Y = 80 else
"111111111111" when X = 126 AND Y = 80 else
"111111111111" when X = 127 AND Y = 80 else
"111111111111" when X = 128 AND Y = 80 else
"111111111111" when X = 129 AND Y = 80 else
"111111111111" when X = 130 AND Y = 80 else
"111111111111" when X = 131 AND Y = 80 else
"111111111111" when X = 132 AND Y = 80 else
"111111111111" when X = 133 AND Y = 80 else
"111111111111" when X = 134 AND Y = 80 else
"111111111111" when X = 135 AND Y = 80 else
"111111111111" when X = 136 AND Y = 80 else
"111111111111" when X = 137 AND Y = 80 else
"111111111111" when X = 138 AND Y = 80 else
"111111111111" when X = 139 AND Y = 80 else
"111111111111" when X = 140 AND Y = 80 else
"111111111111" when X = 141 AND Y = 80 else
"111111111111" when X = 142 AND Y = 80 else
"111111111111" when X = 143 AND Y = 80 else
"111111111111" when X = 144 AND Y = 80 else
"111111111111" when X = 145 AND Y = 80 else
"111111111111" when X = 146 AND Y = 80 else
"111111111111" when X = 147 AND Y = 80 else
"111111111111" when X = 148 AND Y = 80 else
"111111111111" when X = 149 AND Y = 80 else
"111111111111" when X = 150 AND Y = 80 else
"111111111111" when X = 151 AND Y = 80 else
"111111111111" when X = 152 AND Y = 80 else
"111111111111" when X = 153 AND Y = 80 else
"111111111111" when X = 154 AND Y = 80 else
"111111111111" when X = 155 AND Y = 80 else
"111111111111" when X = 156 AND Y = 80 else
"111111111111" when X = 157 AND Y = 80 else
"111111111111" when X = 158 AND Y = 80 else
"111111111111" when X = 159 AND Y = 80 else
"111111111111" when X = 160 AND Y = 80 else
"111111111111" when X = 161 AND Y = 80 else
"111111111111" when X = 162 AND Y = 80 else
"111111111111" when X = 163 AND Y = 80 else
"111111111111" when X = 164 AND Y = 80 else
"111111111111" when X = 165 AND Y = 80 else
"111111111111" when X = 166 AND Y = 80 else
"111111111111" when X = 167 AND Y = 80 else
"111111111111" when X = 168 AND Y = 80 else
"111111111111" when X = 169 AND Y = 80 else
"111111111111" when X = 170 AND Y = 80 else
"111111111111" when X = 171 AND Y = 80 else
"111111111111" when X = 172 AND Y = 80 else
"111111111111" when X = 173 AND Y = 80 else
"111111111111" when X = 174 AND Y = 80 else
"111111111111" when X = 175 AND Y = 80 else
"111111111111" when X = 176 AND Y = 80 else
"111111111111" when X = 177 AND Y = 80 else
"111111111111" when X = 178 AND Y = 80 else
"111111111111" when X = 179 AND Y = 80 else
"111111111111" when X = 180 AND Y = 80 else
"111111111111" when X = 181 AND Y = 80 else
"111111111111" when X = 182 AND Y = 80 else
"111111111111" when X = 183 AND Y = 80 else
"111111111111" when X = 184 AND Y = 80 else
"111111111111" when X = 185 AND Y = 80 else
"111111111111" when X = 186 AND Y = 80 else
"111111111111" when X = 187 AND Y = 80 else
"111111111111" when X = 188 AND Y = 80 else
"111111111111" when X = 189 AND Y = 80 else
"111111111111" when X = 190 AND Y = 80 else
"111111111111" when X = 191 AND Y = 80 else
"111111111111" when X = 192 AND Y = 80 else
"111111111111" when X = 193 AND Y = 80 else
"111111111111" when X = 194 AND Y = 80 else
"111111111111" when X = 195 AND Y = 80 else
"111111111111" when X = 196 AND Y = 80 else
"111111111111" when X = 197 AND Y = 80 else
"111111111111" when X = 198 AND Y = 80 else
"111111111111" when X = 199 AND Y = 80 else
"111111111111" when X = 200 AND Y = 80 else
"111111111111" when X = 201 AND Y = 80 else
"111111111111" when X = 202 AND Y = 80 else
"111111111111" when X = 203 AND Y = 80 else
"111111111111" when X = 204 AND Y = 80 else
"111111111111" when X = 205 AND Y = 80 else
"111111111111" when X = 206 AND Y = 80 else
"111111111111" when X = 207 AND Y = 80 else
"111111111111" when X = 208 AND Y = 80 else
"111111111111" when X = 209 AND Y = 80 else
"111111111111" when X = 210 AND Y = 80 else
"111111111111" when X = 211 AND Y = 80 else
"111111111111" when X = 212 AND Y = 80 else
"111111111111" when X = 213 AND Y = 80 else
"111111111111" when X = 214 AND Y = 80 else
"111111111111" when X = 215 AND Y = 80 else
"111111111111" when X = 216 AND Y = 80 else
"111111111111" when X = 217 AND Y = 80 else
"111111111111" when X = 218 AND Y = 80 else
"111111111111" when X = 219 AND Y = 80 else
"111111111111" when X = 220 AND Y = 80 else
"111111111111" when X = 221 AND Y = 80 else
"111111111111" when X = 222 AND Y = 80 else
"111111111111" when X = 223 AND Y = 80 else
"111111111111" when X = 224 AND Y = 80 else
"111111111111" when X = 225 AND Y = 80 else
"111111111111" when X = 226 AND Y = 80 else
"111111111111" when X = 227 AND Y = 80 else
"111111111111" when X = 228 AND Y = 80 else
"111111111111" when X = 229 AND Y = 80 else
"111111111111" when X = 230 AND Y = 80 else
"111111111111" when X = 231 AND Y = 80 else
"111111111111" when X = 232 AND Y = 80 else
"111111111111" when X = 233 AND Y = 80 else
"111111111111" when X = 234 AND Y = 80 else
"111111111111" when X = 235 AND Y = 80 else
"111111111111" when X = 236 AND Y = 80 else
"111111111111" when X = 237 AND Y = 80 else
"111111111111" when X = 238 AND Y = 80 else
"111111111111" when X = 239 AND Y = 80 else
"111111111111" when X = 240 AND Y = 80 else
"111111111111" when X = 241 AND Y = 80 else
"111111111111" when X = 242 AND Y = 80 else
"111111111111" when X = 243 AND Y = 80 else
"111111111111" when X = 244 AND Y = 80 else
"111111111111" when X = 245 AND Y = 80 else
"111111111111" when X = 246 AND Y = 80 else
"111111111111" when X = 247 AND Y = 80 else
"111111111111" when X = 248 AND Y = 80 else
"111111111111" when X = 249 AND Y = 80 else
"111111111111" when X = 250 AND Y = 80 else
"111111111111" when X = 251 AND Y = 80 else
"111111111111" when X = 252 AND Y = 80 else
"111111111111" when X = 253 AND Y = 80 else
"111111111111" when X = 254 AND Y = 80 else
"111111111111" when X = 255 AND Y = 80 else
"111111111111" when X = 256 AND Y = 80 else
"111111111111" when X = 257 AND Y = 80 else
"111111111111" when X = 258 AND Y = 80 else
"111111111111" when X = 259 AND Y = 80 else
"111111111111" when X = 260 AND Y = 80 else
"111111111111" when X = 261 AND Y = 80 else
"111111111111" when X = 262 AND Y = 80 else
"111111111111" when X = 263 AND Y = 80 else
"111111111111" when X = 264 AND Y = 80 else
"111111111111" when X = 265 AND Y = 80 else
"111111111111" when X = 266 AND Y = 80 else
"111111111111" when X = 267 AND Y = 80 else
"111111111111" when X = 268 AND Y = 80 else
"111111111111" when X = 269 AND Y = 80 else
"110111011111" when X = 270 AND Y = 80 else
"110111011111" when X = 271 AND Y = 80 else
"110111011111" when X = 272 AND Y = 80 else
"110111011111" when X = 273 AND Y = 80 else
"110111011111" when X = 274 AND Y = 80 else
"110111011111" when X = 275 AND Y = 80 else
"110111011111" when X = 276 AND Y = 80 else
"110111011111" when X = 277 AND Y = 80 else
"110111011111" when X = 278 AND Y = 80 else
"110111011111" when X = 279 AND Y = 80 else
"110111011111" when X = 280 AND Y = 80 else
"110111011111" when X = 281 AND Y = 80 else
"110111011111" when X = 282 AND Y = 80 else
"110111011111" when X = 283 AND Y = 80 else
"110111011111" when X = 284 AND Y = 80 else
"110111011111" when X = 285 AND Y = 80 else
"110111011111" when X = 286 AND Y = 80 else
"110111011111" when X = 287 AND Y = 80 else
"110111011111" when X = 288 AND Y = 80 else
"110111011111" when X = 289 AND Y = 80 else
"110111011111" when X = 290 AND Y = 80 else
"110111011111" when X = 291 AND Y = 80 else
"110111011111" when X = 292 AND Y = 80 else
"110111011111" when X = 293 AND Y = 80 else
"110111011111" when X = 294 AND Y = 80 else
"110111011111" when X = 295 AND Y = 80 else
"110111011111" when X = 296 AND Y = 80 else
"110111011111" when X = 297 AND Y = 80 else
"110111011111" when X = 298 AND Y = 80 else
"110111011111" when X = 299 AND Y = 80 else
"110111011111" when X = 300 AND Y = 80 else
"110111011111" when X = 301 AND Y = 80 else
"110111011111" when X = 302 AND Y = 80 else
"110111011111" when X = 303 AND Y = 80 else
"110111011111" when X = 304 AND Y = 80 else
"110111011111" when X = 305 AND Y = 80 else
"110111011111" when X = 306 AND Y = 80 else
"110111011111" when X = 307 AND Y = 80 else
"110111011111" when X = 308 AND Y = 80 else
"110111011111" when X = 309 AND Y = 80 else
"110111011111" when X = 310 AND Y = 80 else
"110111011111" when X = 311 AND Y = 80 else
"110111011111" when X = 312 AND Y = 80 else
"110111011111" when X = 313 AND Y = 80 else
"110111011111" when X = 314 AND Y = 80 else
"110111011111" when X = 315 AND Y = 80 else
"110111011111" when X = 316 AND Y = 80 else
"110111011111" when X = 317 AND Y = 80 else
"110111011111" when X = 318 AND Y = 80 else
"110111011111" when X = 319 AND Y = 80 else
"000000000000" when X = 320 AND Y = 80 else
"000000000000" when X = 321 AND Y = 80 else
"000000000000" when X = 322 AND Y = 80 else
"000000000000" when X = 323 AND Y = 80 else
"000000000000" when X = 324 AND Y = 80 else
"100010011101" when X = 0 AND Y = 81 else
"100010011101" when X = 1 AND Y = 81 else
"100010011101" when X = 2 AND Y = 81 else
"100010011101" when X = 3 AND Y = 81 else
"100010011101" when X = 4 AND Y = 81 else
"100010011101" when X = 5 AND Y = 81 else
"100010011101" when X = 6 AND Y = 81 else
"100010011101" when X = 7 AND Y = 81 else
"100010011101" when X = 8 AND Y = 81 else
"100010011101" when X = 9 AND Y = 81 else
"100010011101" when X = 10 AND Y = 81 else
"100010011101" when X = 11 AND Y = 81 else
"100010011101" when X = 12 AND Y = 81 else
"100010011101" when X = 13 AND Y = 81 else
"100010011101" when X = 14 AND Y = 81 else
"100010011101" when X = 15 AND Y = 81 else
"100010011101" when X = 16 AND Y = 81 else
"100010011101" when X = 17 AND Y = 81 else
"100010011101" when X = 18 AND Y = 81 else
"100010011101" when X = 19 AND Y = 81 else
"100010011101" when X = 20 AND Y = 81 else
"100010011101" when X = 21 AND Y = 81 else
"100010011101" when X = 22 AND Y = 81 else
"100010011101" when X = 23 AND Y = 81 else
"100010011101" when X = 24 AND Y = 81 else
"100010011101" when X = 25 AND Y = 81 else
"100010011101" when X = 26 AND Y = 81 else
"100010011101" when X = 27 AND Y = 81 else
"100010011101" when X = 28 AND Y = 81 else
"100010011101" when X = 29 AND Y = 81 else
"110111011111" when X = 30 AND Y = 81 else
"110111011111" when X = 31 AND Y = 81 else
"110111011111" when X = 32 AND Y = 81 else
"110111011111" when X = 33 AND Y = 81 else
"110111011111" when X = 34 AND Y = 81 else
"110111011111" when X = 35 AND Y = 81 else
"110111011111" when X = 36 AND Y = 81 else
"110111011111" when X = 37 AND Y = 81 else
"110111011111" when X = 38 AND Y = 81 else
"110111011111" when X = 39 AND Y = 81 else
"110111011111" when X = 40 AND Y = 81 else
"110111011111" when X = 41 AND Y = 81 else
"110111011111" when X = 42 AND Y = 81 else
"110111011111" when X = 43 AND Y = 81 else
"110111011111" when X = 44 AND Y = 81 else
"110111011111" when X = 45 AND Y = 81 else
"110111011111" when X = 46 AND Y = 81 else
"110111011111" when X = 47 AND Y = 81 else
"110111011111" when X = 48 AND Y = 81 else
"110111011111" when X = 49 AND Y = 81 else
"110111011111" when X = 50 AND Y = 81 else
"110111011111" when X = 51 AND Y = 81 else
"110111011111" when X = 52 AND Y = 81 else
"110111011111" when X = 53 AND Y = 81 else
"110111011111" when X = 54 AND Y = 81 else
"110111011111" when X = 55 AND Y = 81 else
"110111011111" when X = 56 AND Y = 81 else
"110111011111" when X = 57 AND Y = 81 else
"110111011111" when X = 58 AND Y = 81 else
"110111011111" when X = 59 AND Y = 81 else
"110111011111" when X = 60 AND Y = 81 else
"110111011111" when X = 61 AND Y = 81 else
"110111011111" when X = 62 AND Y = 81 else
"110111011111" when X = 63 AND Y = 81 else
"110111011111" when X = 64 AND Y = 81 else
"110111011111" when X = 65 AND Y = 81 else
"110111011111" when X = 66 AND Y = 81 else
"110111011111" when X = 67 AND Y = 81 else
"110111011111" when X = 68 AND Y = 81 else
"110111011111" when X = 69 AND Y = 81 else
"110111011111" when X = 70 AND Y = 81 else
"110111011111" when X = 71 AND Y = 81 else
"110111011111" when X = 72 AND Y = 81 else
"110111011111" when X = 73 AND Y = 81 else
"110111011111" when X = 74 AND Y = 81 else
"110111011111" when X = 75 AND Y = 81 else
"110111011111" when X = 76 AND Y = 81 else
"110111011111" when X = 77 AND Y = 81 else
"110111011111" when X = 78 AND Y = 81 else
"110111011111" when X = 79 AND Y = 81 else
"110111011111" when X = 80 AND Y = 81 else
"110111011111" when X = 81 AND Y = 81 else
"110111011111" when X = 82 AND Y = 81 else
"110111011111" when X = 83 AND Y = 81 else
"110111011111" when X = 84 AND Y = 81 else
"110111011111" when X = 85 AND Y = 81 else
"110111011111" when X = 86 AND Y = 81 else
"110111011111" when X = 87 AND Y = 81 else
"110111011111" when X = 88 AND Y = 81 else
"110111011111" when X = 89 AND Y = 81 else
"110111011111" when X = 90 AND Y = 81 else
"110111011111" when X = 91 AND Y = 81 else
"110111011111" when X = 92 AND Y = 81 else
"110111011111" when X = 93 AND Y = 81 else
"110111011111" when X = 94 AND Y = 81 else
"110111011111" when X = 95 AND Y = 81 else
"110111011111" when X = 96 AND Y = 81 else
"110111011111" when X = 97 AND Y = 81 else
"110111011111" when X = 98 AND Y = 81 else
"110111011111" when X = 99 AND Y = 81 else
"110111011111" when X = 100 AND Y = 81 else
"110111011111" when X = 101 AND Y = 81 else
"110111011111" when X = 102 AND Y = 81 else
"110111011111" when X = 103 AND Y = 81 else
"110111011111" when X = 104 AND Y = 81 else
"111111111111" when X = 105 AND Y = 81 else
"111111111111" when X = 106 AND Y = 81 else
"111111111111" when X = 107 AND Y = 81 else
"111111111111" when X = 108 AND Y = 81 else
"111111111111" when X = 109 AND Y = 81 else
"111111111111" when X = 110 AND Y = 81 else
"111111111111" when X = 111 AND Y = 81 else
"111111111111" when X = 112 AND Y = 81 else
"111111111111" when X = 113 AND Y = 81 else
"111111111111" when X = 114 AND Y = 81 else
"111111111111" when X = 115 AND Y = 81 else
"111111111111" when X = 116 AND Y = 81 else
"111111111111" when X = 117 AND Y = 81 else
"111111111111" when X = 118 AND Y = 81 else
"111111111111" when X = 119 AND Y = 81 else
"111111111111" when X = 120 AND Y = 81 else
"111111111111" when X = 121 AND Y = 81 else
"111111111111" when X = 122 AND Y = 81 else
"111111111111" when X = 123 AND Y = 81 else
"111111111111" when X = 124 AND Y = 81 else
"111111111111" when X = 125 AND Y = 81 else
"111111111111" when X = 126 AND Y = 81 else
"111111111111" when X = 127 AND Y = 81 else
"111111111111" when X = 128 AND Y = 81 else
"111111111111" when X = 129 AND Y = 81 else
"111111111111" when X = 130 AND Y = 81 else
"111111111111" when X = 131 AND Y = 81 else
"111111111111" when X = 132 AND Y = 81 else
"111111111111" when X = 133 AND Y = 81 else
"111111111111" when X = 134 AND Y = 81 else
"111111111111" when X = 135 AND Y = 81 else
"111111111111" when X = 136 AND Y = 81 else
"111111111111" when X = 137 AND Y = 81 else
"111111111111" when X = 138 AND Y = 81 else
"111111111111" when X = 139 AND Y = 81 else
"111111111111" when X = 140 AND Y = 81 else
"111111111111" when X = 141 AND Y = 81 else
"111111111111" when X = 142 AND Y = 81 else
"111111111111" when X = 143 AND Y = 81 else
"111111111111" when X = 144 AND Y = 81 else
"111111111111" when X = 145 AND Y = 81 else
"111111111111" when X = 146 AND Y = 81 else
"111111111111" when X = 147 AND Y = 81 else
"111111111111" when X = 148 AND Y = 81 else
"111111111111" when X = 149 AND Y = 81 else
"111111111111" when X = 150 AND Y = 81 else
"111111111111" when X = 151 AND Y = 81 else
"111111111111" when X = 152 AND Y = 81 else
"111111111111" when X = 153 AND Y = 81 else
"111111111111" when X = 154 AND Y = 81 else
"111111111111" when X = 155 AND Y = 81 else
"111111111111" when X = 156 AND Y = 81 else
"111111111111" when X = 157 AND Y = 81 else
"111111111111" when X = 158 AND Y = 81 else
"111111111111" when X = 159 AND Y = 81 else
"111111111111" when X = 160 AND Y = 81 else
"111111111111" when X = 161 AND Y = 81 else
"111111111111" when X = 162 AND Y = 81 else
"111111111111" when X = 163 AND Y = 81 else
"111111111111" when X = 164 AND Y = 81 else
"111111111111" when X = 165 AND Y = 81 else
"111111111111" when X = 166 AND Y = 81 else
"111111111111" when X = 167 AND Y = 81 else
"111111111111" when X = 168 AND Y = 81 else
"111111111111" when X = 169 AND Y = 81 else
"111111111111" when X = 170 AND Y = 81 else
"111111111111" when X = 171 AND Y = 81 else
"111111111111" when X = 172 AND Y = 81 else
"111111111111" when X = 173 AND Y = 81 else
"111111111111" when X = 174 AND Y = 81 else
"111111111111" when X = 175 AND Y = 81 else
"111111111111" when X = 176 AND Y = 81 else
"111111111111" when X = 177 AND Y = 81 else
"111111111111" when X = 178 AND Y = 81 else
"111111111111" when X = 179 AND Y = 81 else
"111111111111" when X = 180 AND Y = 81 else
"111111111111" when X = 181 AND Y = 81 else
"111111111111" when X = 182 AND Y = 81 else
"111111111111" when X = 183 AND Y = 81 else
"111111111111" when X = 184 AND Y = 81 else
"111111111111" when X = 185 AND Y = 81 else
"111111111111" when X = 186 AND Y = 81 else
"111111111111" when X = 187 AND Y = 81 else
"111111111111" when X = 188 AND Y = 81 else
"111111111111" when X = 189 AND Y = 81 else
"111111111111" when X = 190 AND Y = 81 else
"111111111111" when X = 191 AND Y = 81 else
"111111111111" when X = 192 AND Y = 81 else
"111111111111" when X = 193 AND Y = 81 else
"111111111111" when X = 194 AND Y = 81 else
"111111111111" when X = 195 AND Y = 81 else
"111111111111" when X = 196 AND Y = 81 else
"111111111111" when X = 197 AND Y = 81 else
"111111111111" when X = 198 AND Y = 81 else
"111111111111" when X = 199 AND Y = 81 else
"111111111111" when X = 200 AND Y = 81 else
"111111111111" when X = 201 AND Y = 81 else
"111111111111" when X = 202 AND Y = 81 else
"111111111111" when X = 203 AND Y = 81 else
"111111111111" when X = 204 AND Y = 81 else
"111111111111" when X = 205 AND Y = 81 else
"111111111111" when X = 206 AND Y = 81 else
"111111111111" when X = 207 AND Y = 81 else
"111111111111" when X = 208 AND Y = 81 else
"111111111111" when X = 209 AND Y = 81 else
"111111111111" when X = 210 AND Y = 81 else
"111111111111" when X = 211 AND Y = 81 else
"111111111111" when X = 212 AND Y = 81 else
"111111111111" when X = 213 AND Y = 81 else
"111111111111" when X = 214 AND Y = 81 else
"111111111111" when X = 215 AND Y = 81 else
"111111111111" when X = 216 AND Y = 81 else
"111111111111" when X = 217 AND Y = 81 else
"111111111111" when X = 218 AND Y = 81 else
"111111111111" when X = 219 AND Y = 81 else
"111111111111" when X = 220 AND Y = 81 else
"111111111111" when X = 221 AND Y = 81 else
"111111111111" when X = 222 AND Y = 81 else
"111111111111" when X = 223 AND Y = 81 else
"111111111111" when X = 224 AND Y = 81 else
"111111111111" when X = 225 AND Y = 81 else
"111111111111" when X = 226 AND Y = 81 else
"111111111111" when X = 227 AND Y = 81 else
"111111111111" when X = 228 AND Y = 81 else
"111111111111" when X = 229 AND Y = 81 else
"111111111111" when X = 230 AND Y = 81 else
"111111111111" when X = 231 AND Y = 81 else
"111111111111" when X = 232 AND Y = 81 else
"111111111111" when X = 233 AND Y = 81 else
"111111111111" when X = 234 AND Y = 81 else
"111111111111" when X = 235 AND Y = 81 else
"111111111111" when X = 236 AND Y = 81 else
"111111111111" when X = 237 AND Y = 81 else
"111111111111" when X = 238 AND Y = 81 else
"111111111111" when X = 239 AND Y = 81 else
"111111111111" when X = 240 AND Y = 81 else
"111111111111" when X = 241 AND Y = 81 else
"111111111111" when X = 242 AND Y = 81 else
"111111111111" when X = 243 AND Y = 81 else
"111111111111" when X = 244 AND Y = 81 else
"111111111111" when X = 245 AND Y = 81 else
"111111111111" when X = 246 AND Y = 81 else
"111111111111" when X = 247 AND Y = 81 else
"111111111111" when X = 248 AND Y = 81 else
"111111111111" when X = 249 AND Y = 81 else
"111111111111" when X = 250 AND Y = 81 else
"111111111111" when X = 251 AND Y = 81 else
"111111111111" when X = 252 AND Y = 81 else
"111111111111" when X = 253 AND Y = 81 else
"111111111111" when X = 254 AND Y = 81 else
"111111111111" when X = 255 AND Y = 81 else
"111111111111" when X = 256 AND Y = 81 else
"111111111111" when X = 257 AND Y = 81 else
"111111111111" when X = 258 AND Y = 81 else
"111111111111" when X = 259 AND Y = 81 else
"111111111111" when X = 260 AND Y = 81 else
"111111111111" when X = 261 AND Y = 81 else
"111111111111" when X = 262 AND Y = 81 else
"111111111111" when X = 263 AND Y = 81 else
"111111111111" when X = 264 AND Y = 81 else
"111111111111" when X = 265 AND Y = 81 else
"111111111111" when X = 266 AND Y = 81 else
"111111111111" when X = 267 AND Y = 81 else
"111111111111" when X = 268 AND Y = 81 else
"111111111111" when X = 269 AND Y = 81 else
"110111011111" when X = 270 AND Y = 81 else
"110111011111" when X = 271 AND Y = 81 else
"110111011111" when X = 272 AND Y = 81 else
"110111011111" when X = 273 AND Y = 81 else
"110111011111" when X = 274 AND Y = 81 else
"110111011111" when X = 275 AND Y = 81 else
"110111011111" when X = 276 AND Y = 81 else
"110111011111" when X = 277 AND Y = 81 else
"110111011111" when X = 278 AND Y = 81 else
"110111011111" when X = 279 AND Y = 81 else
"110111011111" when X = 280 AND Y = 81 else
"110111011111" when X = 281 AND Y = 81 else
"110111011111" when X = 282 AND Y = 81 else
"110111011111" when X = 283 AND Y = 81 else
"110111011111" when X = 284 AND Y = 81 else
"110111011111" when X = 285 AND Y = 81 else
"110111011111" when X = 286 AND Y = 81 else
"110111011111" when X = 287 AND Y = 81 else
"110111011111" when X = 288 AND Y = 81 else
"110111011111" when X = 289 AND Y = 81 else
"110111011111" when X = 290 AND Y = 81 else
"110111011111" when X = 291 AND Y = 81 else
"110111011111" when X = 292 AND Y = 81 else
"110111011111" when X = 293 AND Y = 81 else
"110111011111" when X = 294 AND Y = 81 else
"110111011111" when X = 295 AND Y = 81 else
"110111011111" when X = 296 AND Y = 81 else
"110111011111" when X = 297 AND Y = 81 else
"110111011111" when X = 298 AND Y = 81 else
"110111011111" when X = 299 AND Y = 81 else
"110111011111" when X = 300 AND Y = 81 else
"110111011111" when X = 301 AND Y = 81 else
"110111011111" when X = 302 AND Y = 81 else
"110111011111" when X = 303 AND Y = 81 else
"110111011111" when X = 304 AND Y = 81 else
"110111011111" when X = 305 AND Y = 81 else
"110111011111" when X = 306 AND Y = 81 else
"110111011111" when X = 307 AND Y = 81 else
"110111011111" when X = 308 AND Y = 81 else
"110111011111" when X = 309 AND Y = 81 else
"110111011111" when X = 310 AND Y = 81 else
"110111011111" when X = 311 AND Y = 81 else
"110111011111" when X = 312 AND Y = 81 else
"110111011111" when X = 313 AND Y = 81 else
"110111011111" when X = 314 AND Y = 81 else
"110111011111" when X = 315 AND Y = 81 else
"110111011111" when X = 316 AND Y = 81 else
"110111011111" when X = 317 AND Y = 81 else
"110111011111" when X = 318 AND Y = 81 else
"110111011111" when X = 319 AND Y = 81 else
"000000000000" when X = 320 AND Y = 81 else
"000000000000" when X = 321 AND Y = 81 else
"000000000000" when X = 322 AND Y = 81 else
"000000000000" when X = 323 AND Y = 81 else
"000000000000" when X = 324 AND Y = 81 else
"100010011101" when X = 0 AND Y = 82 else
"100010011101" when X = 1 AND Y = 82 else
"100010011101" when X = 2 AND Y = 82 else
"100010011101" when X = 3 AND Y = 82 else
"100010011101" when X = 4 AND Y = 82 else
"100010011101" when X = 5 AND Y = 82 else
"100010011101" when X = 6 AND Y = 82 else
"100010011101" when X = 7 AND Y = 82 else
"100010011101" when X = 8 AND Y = 82 else
"100010011101" when X = 9 AND Y = 82 else
"100010011101" when X = 10 AND Y = 82 else
"100010011101" when X = 11 AND Y = 82 else
"100010011101" when X = 12 AND Y = 82 else
"100010011101" when X = 13 AND Y = 82 else
"100010011101" when X = 14 AND Y = 82 else
"100010011101" when X = 15 AND Y = 82 else
"100010011101" when X = 16 AND Y = 82 else
"100010011101" when X = 17 AND Y = 82 else
"100010011101" when X = 18 AND Y = 82 else
"100010011101" when X = 19 AND Y = 82 else
"100010011101" when X = 20 AND Y = 82 else
"100010011101" when X = 21 AND Y = 82 else
"100010011101" when X = 22 AND Y = 82 else
"100010011101" when X = 23 AND Y = 82 else
"100010011101" when X = 24 AND Y = 82 else
"100010011101" when X = 25 AND Y = 82 else
"100010011101" when X = 26 AND Y = 82 else
"100010011101" when X = 27 AND Y = 82 else
"100010011101" when X = 28 AND Y = 82 else
"100010011101" when X = 29 AND Y = 82 else
"110111011111" when X = 30 AND Y = 82 else
"110111011111" when X = 31 AND Y = 82 else
"110111011111" when X = 32 AND Y = 82 else
"110111011111" when X = 33 AND Y = 82 else
"110111011111" when X = 34 AND Y = 82 else
"110111011111" when X = 35 AND Y = 82 else
"110111011111" when X = 36 AND Y = 82 else
"110111011111" when X = 37 AND Y = 82 else
"110111011111" when X = 38 AND Y = 82 else
"110111011111" when X = 39 AND Y = 82 else
"110111011111" when X = 40 AND Y = 82 else
"110111011111" when X = 41 AND Y = 82 else
"110111011111" when X = 42 AND Y = 82 else
"110111011111" when X = 43 AND Y = 82 else
"110111011111" when X = 44 AND Y = 82 else
"110111011111" when X = 45 AND Y = 82 else
"110111011111" when X = 46 AND Y = 82 else
"110111011111" when X = 47 AND Y = 82 else
"110111011111" when X = 48 AND Y = 82 else
"110111011111" when X = 49 AND Y = 82 else
"110111011111" when X = 50 AND Y = 82 else
"110111011111" when X = 51 AND Y = 82 else
"110111011111" when X = 52 AND Y = 82 else
"110111011111" when X = 53 AND Y = 82 else
"110111011111" when X = 54 AND Y = 82 else
"110111011111" when X = 55 AND Y = 82 else
"110111011111" when X = 56 AND Y = 82 else
"110111011111" when X = 57 AND Y = 82 else
"110111011111" when X = 58 AND Y = 82 else
"110111011111" when X = 59 AND Y = 82 else
"110111011111" when X = 60 AND Y = 82 else
"110111011111" when X = 61 AND Y = 82 else
"110111011111" when X = 62 AND Y = 82 else
"110111011111" when X = 63 AND Y = 82 else
"110111011111" when X = 64 AND Y = 82 else
"110111011111" when X = 65 AND Y = 82 else
"110111011111" when X = 66 AND Y = 82 else
"110111011111" when X = 67 AND Y = 82 else
"110111011111" when X = 68 AND Y = 82 else
"110111011111" when X = 69 AND Y = 82 else
"110111011111" when X = 70 AND Y = 82 else
"110111011111" when X = 71 AND Y = 82 else
"110111011111" when X = 72 AND Y = 82 else
"110111011111" when X = 73 AND Y = 82 else
"110111011111" when X = 74 AND Y = 82 else
"110111011111" when X = 75 AND Y = 82 else
"110111011111" when X = 76 AND Y = 82 else
"110111011111" when X = 77 AND Y = 82 else
"110111011111" when X = 78 AND Y = 82 else
"110111011111" when X = 79 AND Y = 82 else
"110111011111" when X = 80 AND Y = 82 else
"110111011111" when X = 81 AND Y = 82 else
"110111011111" when X = 82 AND Y = 82 else
"110111011111" when X = 83 AND Y = 82 else
"110111011111" when X = 84 AND Y = 82 else
"110111011111" when X = 85 AND Y = 82 else
"110111011111" when X = 86 AND Y = 82 else
"110111011111" when X = 87 AND Y = 82 else
"110111011111" when X = 88 AND Y = 82 else
"110111011111" when X = 89 AND Y = 82 else
"110111011111" when X = 90 AND Y = 82 else
"110111011111" when X = 91 AND Y = 82 else
"110111011111" when X = 92 AND Y = 82 else
"110111011111" when X = 93 AND Y = 82 else
"110111011111" when X = 94 AND Y = 82 else
"110111011111" when X = 95 AND Y = 82 else
"110111011111" when X = 96 AND Y = 82 else
"110111011111" when X = 97 AND Y = 82 else
"110111011111" when X = 98 AND Y = 82 else
"110111011111" when X = 99 AND Y = 82 else
"110111011111" when X = 100 AND Y = 82 else
"110111011111" when X = 101 AND Y = 82 else
"110111011111" when X = 102 AND Y = 82 else
"110111011111" when X = 103 AND Y = 82 else
"110111011111" when X = 104 AND Y = 82 else
"111111111111" when X = 105 AND Y = 82 else
"111111111111" when X = 106 AND Y = 82 else
"111111111111" when X = 107 AND Y = 82 else
"111111111111" when X = 108 AND Y = 82 else
"111111111111" when X = 109 AND Y = 82 else
"111111111111" when X = 110 AND Y = 82 else
"111111111111" when X = 111 AND Y = 82 else
"111111111111" when X = 112 AND Y = 82 else
"111111111111" when X = 113 AND Y = 82 else
"111111111111" when X = 114 AND Y = 82 else
"111111111111" when X = 115 AND Y = 82 else
"111111111111" when X = 116 AND Y = 82 else
"111111111111" when X = 117 AND Y = 82 else
"111111111111" when X = 118 AND Y = 82 else
"111111111111" when X = 119 AND Y = 82 else
"111111111111" when X = 120 AND Y = 82 else
"111111111111" when X = 121 AND Y = 82 else
"111111111111" when X = 122 AND Y = 82 else
"111111111111" when X = 123 AND Y = 82 else
"111111111111" when X = 124 AND Y = 82 else
"111111111111" when X = 125 AND Y = 82 else
"111111111111" when X = 126 AND Y = 82 else
"111111111111" when X = 127 AND Y = 82 else
"111111111111" when X = 128 AND Y = 82 else
"111111111111" when X = 129 AND Y = 82 else
"111111111111" when X = 130 AND Y = 82 else
"111111111111" when X = 131 AND Y = 82 else
"111111111111" when X = 132 AND Y = 82 else
"111111111111" when X = 133 AND Y = 82 else
"111111111111" when X = 134 AND Y = 82 else
"111111111111" when X = 135 AND Y = 82 else
"111111111111" when X = 136 AND Y = 82 else
"111111111111" when X = 137 AND Y = 82 else
"111111111111" when X = 138 AND Y = 82 else
"111111111111" when X = 139 AND Y = 82 else
"111111111111" when X = 140 AND Y = 82 else
"111111111111" when X = 141 AND Y = 82 else
"111111111111" when X = 142 AND Y = 82 else
"111111111111" when X = 143 AND Y = 82 else
"111111111111" when X = 144 AND Y = 82 else
"111111111111" when X = 145 AND Y = 82 else
"111111111111" when X = 146 AND Y = 82 else
"111111111111" when X = 147 AND Y = 82 else
"111111111111" when X = 148 AND Y = 82 else
"111111111111" when X = 149 AND Y = 82 else
"111111111111" when X = 150 AND Y = 82 else
"111111111111" when X = 151 AND Y = 82 else
"111111111111" when X = 152 AND Y = 82 else
"111111111111" when X = 153 AND Y = 82 else
"111111111111" when X = 154 AND Y = 82 else
"111111111111" when X = 155 AND Y = 82 else
"111111111111" when X = 156 AND Y = 82 else
"111111111111" when X = 157 AND Y = 82 else
"111111111111" when X = 158 AND Y = 82 else
"111111111111" when X = 159 AND Y = 82 else
"111111111111" when X = 160 AND Y = 82 else
"111111111111" when X = 161 AND Y = 82 else
"111111111111" when X = 162 AND Y = 82 else
"111111111111" when X = 163 AND Y = 82 else
"111111111111" when X = 164 AND Y = 82 else
"111111111111" when X = 165 AND Y = 82 else
"111111111111" when X = 166 AND Y = 82 else
"111111111111" when X = 167 AND Y = 82 else
"111111111111" when X = 168 AND Y = 82 else
"111111111111" when X = 169 AND Y = 82 else
"111111111111" when X = 170 AND Y = 82 else
"111111111111" when X = 171 AND Y = 82 else
"111111111111" when X = 172 AND Y = 82 else
"111111111111" when X = 173 AND Y = 82 else
"111111111111" when X = 174 AND Y = 82 else
"111111111111" when X = 175 AND Y = 82 else
"111111111111" when X = 176 AND Y = 82 else
"111111111111" when X = 177 AND Y = 82 else
"111111111111" when X = 178 AND Y = 82 else
"111111111111" when X = 179 AND Y = 82 else
"111111111111" when X = 180 AND Y = 82 else
"111111111111" when X = 181 AND Y = 82 else
"111111111111" when X = 182 AND Y = 82 else
"111111111111" when X = 183 AND Y = 82 else
"111111111111" when X = 184 AND Y = 82 else
"111111111111" when X = 185 AND Y = 82 else
"111111111111" when X = 186 AND Y = 82 else
"111111111111" when X = 187 AND Y = 82 else
"111111111111" when X = 188 AND Y = 82 else
"111111111111" when X = 189 AND Y = 82 else
"111111111111" when X = 190 AND Y = 82 else
"111111111111" when X = 191 AND Y = 82 else
"111111111111" when X = 192 AND Y = 82 else
"111111111111" when X = 193 AND Y = 82 else
"111111111111" when X = 194 AND Y = 82 else
"111111111111" when X = 195 AND Y = 82 else
"111111111111" when X = 196 AND Y = 82 else
"111111111111" when X = 197 AND Y = 82 else
"111111111111" when X = 198 AND Y = 82 else
"111111111111" when X = 199 AND Y = 82 else
"111111111111" when X = 200 AND Y = 82 else
"111111111111" when X = 201 AND Y = 82 else
"111111111111" when X = 202 AND Y = 82 else
"111111111111" when X = 203 AND Y = 82 else
"111111111111" when X = 204 AND Y = 82 else
"111111111111" when X = 205 AND Y = 82 else
"111111111111" when X = 206 AND Y = 82 else
"111111111111" when X = 207 AND Y = 82 else
"111111111111" when X = 208 AND Y = 82 else
"111111111111" when X = 209 AND Y = 82 else
"111111111111" when X = 210 AND Y = 82 else
"111111111111" when X = 211 AND Y = 82 else
"111111111111" when X = 212 AND Y = 82 else
"111111111111" when X = 213 AND Y = 82 else
"111111111111" when X = 214 AND Y = 82 else
"111111111111" when X = 215 AND Y = 82 else
"111111111111" when X = 216 AND Y = 82 else
"111111111111" when X = 217 AND Y = 82 else
"111111111111" when X = 218 AND Y = 82 else
"111111111111" when X = 219 AND Y = 82 else
"111111111111" when X = 220 AND Y = 82 else
"111111111111" when X = 221 AND Y = 82 else
"111111111111" when X = 222 AND Y = 82 else
"111111111111" when X = 223 AND Y = 82 else
"111111111111" when X = 224 AND Y = 82 else
"111111111111" when X = 225 AND Y = 82 else
"111111111111" when X = 226 AND Y = 82 else
"111111111111" when X = 227 AND Y = 82 else
"111111111111" when X = 228 AND Y = 82 else
"111111111111" when X = 229 AND Y = 82 else
"111111111111" when X = 230 AND Y = 82 else
"111111111111" when X = 231 AND Y = 82 else
"111111111111" when X = 232 AND Y = 82 else
"111111111111" when X = 233 AND Y = 82 else
"111111111111" when X = 234 AND Y = 82 else
"111111111111" when X = 235 AND Y = 82 else
"111111111111" when X = 236 AND Y = 82 else
"111111111111" when X = 237 AND Y = 82 else
"111111111111" when X = 238 AND Y = 82 else
"111111111111" when X = 239 AND Y = 82 else
"111111111111" when X = 240 AND Y = 82 else
"111111111111" when X = 241 AND Y = 82 else
"111111111111" when X = 242 AND Y = 82 else
"111111111111" when X = 243 AND Y = 82 else
"111111111111" when X = 244 AND Y = 82 else
"111111111111" when X = 245 AND Y = 82 else
"111111111111" when X = 246 AND Y = 82 else
"111111111111" when X = 247 AND Y = 82 else
"111111111111" when X = 248 AND Y = 82 else
"111111111111" when X = 249 AND Y = 82 else
"111111111111" when X = 250 AND Y = 82 else
"111111111111" when X = 251 AND Y = 82 else
"111111111111" when X = 252 AND Y = 82 else
"111111111111" when X = 253 AND Y = 82 else
"111111111111" when X = 254 AND Y = 82 else
"111111111111" when X = 255 AND Y = 82 else
"111111111111" when X = 256 AND Y = 82 else
"111111111111" when X = 257 AND Y = 82 else
"111111111111" when X = 258 AND Y = 82 else
"111111111111" when X = 259 AND Y = 82 else
"111111111111" when X = 260 AND Y = 82 else
"111111111111" when X = 261 AND Y = 82 else
"111111111111" when X = 262 AND Y = 82 else
"111111111111" when X = 263 AND Y = 82 else
"111111111111" when X = 264 AND Y = 82 else
"111111111111" when X = 265 AND Y = 82 else
"111111111111" when X = 266 AND Y = 82 else
"111111111111" when X = 267 AND Y = 82 else
"111111111111" when X = 268 AND Y = 82 else
"111111111111" when X = 269 AND Y = 82 else
"110111011111" when X = 270 AND Y = 82 else
"110111011111" when X = 271 AND Y = 82 else
"110111011111" when X = 272 AND Y = 82 else
"110111011111" when X = 273 AND Y = 82 else
"110111011111" when X = 274 AND Y = 82 else
"110111011111" when X = 275 AND Y = 82 else
"110111011111" when X = 276 AND Y = 82 else
"110111011111" when X = 277 AND Y = 82 else
"110111011111" when X = 278 AND Y = 82 else
"110111011111" when X = 279 AND Y = 82 else
"110111011111" when X = 280 AND Y = 82 else
"110111011111" when X = 281 AND Y = 82 else
"110111011111" when X = 282 AND Y = 82 else
"110111011111" when X = 283 AND Y = 82 else
"110111011111" when X = 284 AND Y = 82 else
"110111011111" when X = 285 AND Y = 82 else
"110111011111" when X = 286 AND Y = 82 else
"110111011111" when X = 287 AND Y = 82 else
"110111011111" when X = 288 AND Y = 82 else
"110111011111" when X = 289 AND Y = 82 else
"110111011111" when X = 290 AND Y = 82 else
"110111011111" when X = 291 AND Y = 82 else
"110111011111" when X = 292 AND Y = 82 else
"110111011111" when X = 293 AND Y = 82 else
"110111011111" when X = 294 AND Y = 82 else
"110111011111" when X = 295 AND Y = 82 else
"110111011111" when X = 296 AND Y = 82 else
"110111011111" when X = 297 AND Y = 82 else
"110111011111" when X = 298 AND Y = 82 else
"110111011111" when X = 299 AND Y = 82 else
"110111011111" when X = 300 AND Y = 82 else
"110111011111" when X = 301 AND Y = 82 else
"110111011111" when X = 302 AND Y = 82 else
"110111011111" when X = 303 AND Y = 82 else
"110111011111" when X = 304 AND Y = 82 else
"110111011111" when X = 305 AND Y = 82 else
"110111011111" when X = 306 AND Y = 82 else
"110111011111" when X = 307 AND Y = 82 else
"110111011111" when X = 308 AND Y = 82 else
"110111011111" when X = 309 AND Y = 82 else
"110111011111" when X = 310 AND Y = 82 else
"110111011111" when X = 311 AND Y = 82 else
"110111011111" when X = 312 AND Y = 82 else
"110111011111" when X = 313 AND Y = 82 else
"110111011111" when X = 314 AND Y = 82 else
"110111011111" when X = 315 AND Y = 82 else
"110111011111" when X = 316 AND Y = 82 else
"110111011111" when X = 317 AND Y = 82 else
"110111011111" when X = 318 AND Y = 82 else
"110111011111" when X = 319 AND Y = 82 else
"000000000000" when X = 320 AND Y = 82 else
"000000000000" when X = 321 AND Y = 82 else
"000000000000" when X = 322 AND Y = 82 else
"000000000000" when X = 323 AND Y = 82 else
"000000000000" when X = 324 AND Y = 82 else
"100010011101" when X = 0 AND Y = 83 else
"100010011101" when X = 1 AND Y = 83 else
"100010011101" when X = 2 AND Y = 83 else
"100010011101" when X = 3 AND Y = 83 else
"100010011101" when X = 4 AND Y = 83 else
"100010011101" when X = 5 AND Y = 83 else
"100010011101" when X = 6 AND Y = 83 else
"100010011101" when X = 7 AND Y = 83 else
"100010011101" when X = 8 AND Y = 83 else
"100010011101" when X = 9 AND Y = 83 else
"100010011101" when X = 10 AND Y = 83 else
"100010011101" when X = 11 AND Y = 83 else
"100010011101" when X = 12 AND Y = 83 else
"100010011101" when X = 13 AND Y = 83 else
"100010011101" when X = 14 AND Y = 83 else
"100010011101" when X = 15 AND Y = 83 else
"100010011101" when X = 16 AND Y = 83 else
"100010011101" when X = 17 AND Y = 83 else
"100010011101" when X = 18 AND Y = 83 else
"100010011101" when X = 19 AND Y = 83 else
"100010011101" when X = 20 AND Y = 83 else
"100010011101" when X = 21 AND Y = 83 else
"100010011101" when X = 22 AND Y = 83 else
"100010011101" when X = 23 AND Y = 83 else
"100010011101" when X = 24 AND Y = 83 else
"100010011101" when X = 25 AND Y = 83 else
"100010011101" when X = 26 AND Y = 83 else
"100010011101" when X = 27 AND Y = 83 else
"100010011101" when X = 28 AND Y = 83 else
"100010011101" when X = 29 AND Y = 83 else
"110111011111" when X = 30 AND Y = 83 else
"110111011111" when X = 31 AND Y = 83 else
"110111011111" when X = 32 AND Y = 83 else
"110111011111" when X = 33 AND Y = 83 else
"110111011111" when X = 34 AND Y = 83 else
"110111011111" when X = 35 AND Y = 83 else
"110111011111" when X = 36 AND Y = 83 else
"110111011111" when X = 37 AND Y = 83 else
"110111011111" when X = 38 AND Y = 83 else
"110111011111" when X = 39 AND Y = 83 else
"110111011111" when X = 40 AND Y = 83 else
"110111011111" when X = 41 AND Y = 83 else
"110111011111" when X = 42 AND Y = 83 else
"110111011111" when X = 43 AND Y = 83 else
"110111011111" when X = 44 AND Y = 83 else
"110111011111" when X = 45 AND Y = 83 else
"110111011111" when X = 46 AND Y = 83 else
"110111011111" when X = 47 AND Y = 83 else
"110111011111" when X = 48 AND Y = 83 else
"110111011111" when X = 49 AND Y = 83 else
"110111011111" when X = 50 AND Y = 83 else
"110111011111" when X = 51 AND Y = 83 else
"110111011111" when X = 52 AND Y = 83 else
"110111011111" when X = 53 AND Y = 83 else
"110111011111" when X = 54 AND Y = 83 else
"110111011111" when X = 55 AND Y = 83 else
"110111011111" when X = 56 AND Y = 83 else
"110111011111" when X = 57 AND Y = 83 else
"110111011111" when X = 58 AND Y = 83 else
"110111011111" when X = 59 AND Y = 83 else
"110111011111" when X = 60 AND Y = 83 else
"110111011111" when X = 61 AND Y = 83 else
"110111011111" when X = 62 AND Y = 83 else
"110111011111" when X = 63 AND Y = 83 else
"110111011111" when X = 64 AND Y = 83 else
"110111011111" when X = 65 AND Y = 83 else
"110111011111" when X = 66 AND Y = 83 else
"110111011111" when X = 67 AND Y = 83 else
"110111011111" when X = 68 AND Y = 83 else
"110111011111" when X = 69 AND Y = 83 else
"110111011111" when X = 70 AND Y = 83 else
"110111011111" when X = 71 AND Y = 83 else
"110111011111" when X = 72 AND Y = 83 else
"110111011111" when X = 73 AND Y = 83 else
"110111011111" when X = 74 AND Y = 83 else
"110111011111" when X = 75 AND Y = 83 else
"110111011111" when X = 76 AND Y = 83 else
"110111011111" when X = 77 AND Y = 83 else
"110111011111" when X = 78 AND Y = 83 else
"110111011111" when X = 79 AND Y = 83 else
"110111011111" when X = 80 AND Y = 83 else
"110111011111" when X = 81 AND Y = 83 else
"110111011111" when X = 82 AND Y = 83 else
"110111011111" when X = 83 AND Y = 83 else
"110111011111" when X = 84 AND Y = 83 else
"110111011111" when X = 85 AND Y = 83 else
"110111011111" when X = 86 AND Y = 83 else
"110111011111" when X = 87 AND Y = 83 else
"110111011111" when X = 88 AND Y = 83 else
"110111011111" when X = 89 AND Y = 83 else
"110111011111" when X = 90 AND Y = 83 else
"110111011111" when X = 91 AND Y = 83 else
"110111011111" when X = 92 AND Y = 83 else
"110111011111" when X = 93 AND Y = 83 else
"110111011111" when X = 94 AND Y = 83 else
"110111011111" when X = 95 AND Y = 83 else
"110111011111" when X = 96 AND Y = 83 else
"110111011111" when X = 97 AND Y = 83 else
"110111011111" when X = 98 AND Y = 83 else
"110111011111" when X = 99 AND Y = 83 else
"110111011111" when X = 100 AND Y = 83 else
"110111011111" when X = 101 AND Y = 83 else
"110111011111" when X = 102 AND Y = 83 else
"110111011111" when X = 103 AND Y = 83 else
"110111011111" when X = 104 AND Y = 83 else
"111111111111" when X = 105 AND Y = 83 else
"111111111111" when X = 106 AND Y = 83 else
"111111111111" when X = 107 AND Y = 83 else
"111111111111" when X = 108 AND Y = 83 else
"111111111111" when X = 109 AND Y = 83 else
"111111111111" when X = 110 AND Y = 83 else
"111111111111" when X = 111 AND Y = 83 else
"111111111111" when X = 112 AND Y = 83 else
"111111111111" when X = 113 AND Y = 83 else
"111111111111" when X = 114 AND Y = 83 else
"111111111111" when X = 115 AND Y = 83 else
"111111111111" when X = 116 AND Y = 83 else
"111111111111" when X = 117 AND Y = 83 else
"111111111111" when X = 118 AND Y = 83 else
"111111111111" when X = 119 AND Y = 83 else
"111111111111" when X = 120 AND Y = 83 else
"111111111111" when X = 121 AND Y = 83 else
"111111111111" when X = 122 AND Y = 83 else
"111111111111" when X = 123 AND Y = 83 else
"111111111111" when X = 124 AND Y = 83 else
"111111111111" when X = 125 AND Y = 83 else
"111111111111" when X = 126 AND Y = 83 else
"111111111111" when X = 127 AND Y = 83 else
"111111111111" when X = 128 AND Y = 83 else
"111111111111" when X = 129 AND Y = 83 else
"111111111111" when X = 130 AND Y = 83 else
"111111111111" when X = 131 AND Y = 83 else
"111111111111" when X = 132 AND Y = 83 else
"111111111111" when X = 133 AND Y = 83 else
"111111111111" when X = 134 AND Y = 83 else
"111111111111" when X = 135 AND Y = 83 else
"111111111111" when X = 136 AND Y = 83 else
"111111111111" when X = 137 AND Y = 83 else
"111111111111" when X = 138 AND Y = 83 else
"111111111111" when X = 139 AND Y = 83 else
"111111111111" when X = 140 AND Y = 83 else
"111111111111" when X = 141 AND Y = 83 else
"111111111111" when X = 142 AND Y = 83 else
"111111111111" when X = 143 AND Y = 83 else
"111111111111" when X = 144 AND Y = 83 else
"111111111111" when X = 145 AND Y = 83 else
"111111111111" when X = 146 AND Y = 83 else
"111111111111" when X = 147 AND Y = 83 else
"111111111111" when X = 148 AND Y = 83 else
"111111111111" when X = 149 AND Y = 83 else
"111111111111" when X = 150 AND Y = 83 else
"111111111111" when X = 151 AND Y = 83 else
"111111111111" when X = 152 AND Y = 83 else
"111111111111" when X = 153 AND Y = 83 else
"111111111111" when X = 154 AND Y = 83 else
"111111111111" when X = 155 AND Y = 83 else
"111111111111" when X = 156 AND Y = 83 else
"111111111111" when X = 157 AND Y = 83 else
"111111111111" when X = 158 AND Y = 83 else
"111111111111" when X = 159 AND Y = 83 else
"111111111111" when X = 160 AND Y = 83 else
"111111111111" when X = 161 AND Y = 83 else
"111111111111" when X = 162 AND Y = 83 else
"111111111111" when X = 163 AND Y = 83 else
"111111111111" when X = 164 AND Y = 83 else
"111111111111" when X = 165 AND Y = 83 else
"111111111111" when X = 166 AND Y = 83 else
"111111111111" when X = 167 AND Y = 83 else
"111111111111" when X = 168 AND Y = 83 else
"111111111111" when X = 169 AND Y = 83 else
"111111111111" when X = 170 AND Y = 83 else
"111111111111" when X = 171 AND Y = 83 else
"111111111111" when X = 172 AND Y = 83 else
"111111111111" when X = 173 AND Y = 83 else
"111111111111" when X = 174 AND Y = 83 else
"111111111111" when X = 175 AND Y = 83 else
"111111111111" when X = 176 AND Y = 83 else
"111111111111" when X = 177 AND Y = 83 else
"111111111111" when X = 178 AND Y = 83 else
"111111111111" when X = 179 AND Y = 83 else
"111111111111" when X = 180 AND Y = 83 else
"111111111111" when X = 181 AND Y = 83 else
"111111111111" when X = 182 AND Y = 83 else
"111111111111" when X = 183 AND Y = 83 else
"111111111111" when X = 184 AND Y = 83 else
"111111111111" when X = 185 AND Y = 83 else
"111111111111" when X = 186 AND Y = 83 else
"111111111111" when X = 187 AND Y = 83 else
"111111111111" when X = 188 AND Y = 83 else
"111111111111" when X = 189 AND Y = 83 else
"111111111111" when X = 190 AND Y = 83 else
"111111111111" when X = 191 AND Y = 83 else
"111111111111" when X = 192 AND Y = 83 else
"111111111111" when X = 193 AND Y = 83 else
"111111111111" when X = 194 AND Y = 83 else
"111111111111" when X = 195 AND Y = 83 else
"111111111111" when X = 196 AND Y = 83 else
"111111111111" when X = 197 AND Y = 83 else
"111111111111" when X = 198 AND Y = 83 else
"111111111111" when X = 199 AND Y = 83 else
"111111111111" when X = 200 AND Y = 83 else
"111111111111" when X = 201 AND Y = 83 else
"111111111111" when X = 202 AND Y = 83 else
"111111111111" when X = 203 AND Y = 83 else
"111111111111" when X = 204 AND Y = 83 else
"111111111111" when X = 205 AND Y = 83 else
"111111111111" when X = 206 AND Y = 83 else
"111111111111" when X = 207 AND Y = 83 else
"111111111111" when X = 208 AND Y = 83 else
"111111111111" when X = 209 AND Y = 83 else
"111111111111" when X = 210 AND Y = 83 else
"111111111111" when X = 211 AND Y = 83 else
"111111111111" when X = 212 AND Y = 83 else
"111111111111" when X = 213 AND Y = 83 else
"111111111111" when X = 214 AND Y = 83 else
"111111111111" when X = 215 AND Y = 83 else
"111111111111" when X = 216 AND Y = 83 else
"111111111111" when X = 217 AND Y = 83 else
"111111111111" when X = 218 AND Y = 83 else
"111111111111" when X = 219 AND Y = 83 else
"111111111111" when X = 220 AND Y = 83 else
"111111111111" when X = 221 AND Y = 83 else
"111111111111" when X = 222 AND Y = 83 else
"111111111111" when X = 223 AND Y = 83 else
"111111111111" when X = 224 AND Y = 83 else
"111111111111" when X = 225 AND Y = 83 else
"111111111111" when X = 226 AND Y = 83 else
"111111111111" when X = 227 AND Y = 83 else
"111111111111" when X = 228 AND Y = 83 else
"111111111111" when X = 229 AND Y = 83 else
"111111111111" when X = 230 AND Y = 83 else
"111111111111" when X = 231 AND Y = 83 else
"111111111111" when X = 232 AND Y = 83 else
"111111111111" when X = 233 AND Y = 83 else
"111111111111" when X = 234 AND Y = 83 else
"111111111111" when X = 235 AND Y = 83 else
"111111111111" when X = 236 AND Y = 83 else
"111111111111" when X = 237 AND Y = 83 else
"111111111111" when X = 238 AND Y = 83 else
"111111111111" when X = 239 AND Y = 83 else
"111111111111" when X = 240 AND Y = 83 else
"111111111111" when X = 241 AND Y = 83 else
"111111111111" when X = 242 AND Y = 83 else
"111111111111" when X = 243 AND Y = 83 else
"111111111111" when X = 244 AND Y = 83 else
"111111111111" when X = 245 AND Y = 83 else
"111111111111" when X = 246 AND Y = 83 else
"111111111111" when X = 247 AND Y = 83 else
"111111111111" when X = 248 AND Y = 83 else
"111111111111" when X = 249 AND Y = 83 else
"111111111111" when X = 250 AND Y = 83 else
"111111111111" when X = 251 AND Y = 83 else
"111111111111" when X = 252 AND Y = 83 else
"111111111111" when X = 253 AND Y = 83 else
"111111111111" when X = 254 AND Y = 83 else
"111111111111" when X = 255 AND Y = 83 else
"111111111111" when X = 256 AND Y = 83 else
"111111111111" when X = 257 AND Y = 83 else
"111111111111" when X = 258 AND Y = 83 else
"111111111111" when X = 259 AND Y = 83 else
"111111111111" when X = 260 AND Y = 83 else
"111111111111" when X = 261 AND Y = 83 else
"111111111111" when X = 262 AND Y = 83 else
"111111111111" when X = 263 AND Y = 83 else
"111111111111" when X = 264 AND Y = 83 else
"111111111111" when X = 265 AND Y = 83 else
"111111111111" when X = 266 AND Y = 83 else
"111111111111" when X = 267 AND Y = 83 else
"111111111111" when X = 268 AND Y = 83 else
"111111111111" when X = 269 AND Y = 83 else
"110111011111" when X = 270 AND Y = 83 else
"110111011111" when X = 271 AND Y = 83 else
"110111011111" when X = 272 AND Y = 83 else
"110111011111" when X = 273 AND Y = 83 else
"110111011111" when X = 274 AND Y = 83 else
"110111011111" when X = 275 AND Y = 83 else
"110111011111" when X = 276 AND Y = 83 else
"110111011111" when X = 277 AND Y = 83 else
"110111011111" when X = 278 AND Y = 83 else
"110111011111" when X = 279 AND Y = 83 else
"110111011111" when X = 280 AND Y = 83 else
"110111011111" when X = 281 AND Y = 83 else
"110111011111" when X = 282 AND Y = 83 else
"110111011111" when X = 283 AND Y = 83 else
"110111011111" when X = 284 AND Y = 83 else
"110111011111" when X = 285 AND Y = 83 else
"110111011111" when X = 286 AND Y = 83 else
"110111011111" when X = 287 AND Y = 83 else
"110111011111" when X = 288 AND Y = 83 else
"110111011111" when X = 289 AND Y = 83 else
"110111011111" when X = 290 AND Y = 83 else
"110111011111" when X = 291 AND Y = 83 else
"110111011111" when X = 292 AND Y = 83 else
"110111011111" when X = 293 AND Y = 83 else
"110111011111" when X = 294 AND Y = 83 else
"110111011111" when X = 295 AND Y = 83 else
"110111011111" when X = 296 AND Y = 83 else
"110111011111" when X = 297 AND Y = 83 else
"110111011111" when X = 298 AND Y = 83 else
"110111011111" when X = 299 AND Y = 83 else
"110111011111" when X = 300 AND Y = 83 else
"110111011111" when X = 301 AND Y = 83 else
"110111011111" when X = 302 AND Y = 83 else
"110111011111" when X = 303 AND Y = 83 else
"110111011111" when X = 304 AND Y = 83 else
"110111011111" when X = 305 AND Y = 83 else
"110111011111" when X = 306 AND Y = 83 else
"110111011111" when X = 307 AND Y = 83 else
"110111011111" when X = 308 AND Y = 83 else
"110111011111" when X = 309 AND Y = 83 else
"110111011111" when X = 310 AND Y = 83 else
"110111011111" when X = 311 AND Y = 83 else
"110111011111" when X = 312 AND Y = 83 else
"110111011111" when X = 313 AND Y = 83 else
"110111011111" when X = 314 AND Y = 83 else
"110111011111" when X = 315 AND Y = 83 else
"110111011111" when X = 316 AND Y = 83 else
"110111011111" when X = 317 AND Y = 83 else
"110111011111" when X = 318 AND Y = 83 else
"110111011111" when X = 319 AND Y = 83 else
"000000000000" when X = 320 AND Y = 83 else
"000000000000" when X = 321 AND Y = 83 else
"000000000000" when X = 322 AND Y = 83 else
"000000000000" when X = 323 AND Y = 83 else
"000000000000" when X = 324 AND Y = 83 else
"100010011101" when X = 0 AND Y = 84 else
"100010011101" when X = 1 AND Y = 84 else
"100010011101" when X = 2 AND Y = 84 else
"100010011101" when X = 3 AND Y = 84 else
"100010011101" when X = 4 AND Y = 84 else
"100010011101" when X = 5 AND Y = 84 else
"100010011101" when X = 6 AND Y = 84 else
"100010011101" when X = 7 AND Y = 84 else
"100010011101" when X = 8 AND Y = 84 else
"100010011101" when X = 9 AND Y = 84 else
"100010011101" when X = 10 AND Y = 84 else
"100010011101" when X = 11 AND Y = 84 else
"100010011101" when X = 12 AND Y = 84 else
"100010011101" when X = 13 AND Y = 84 else
"100010011101" when X = 14 AND Y = 84 else
"100010011101" when X = 15 AND Y = 84 else
"100010011101" when X = 16 AND Y = 84 else
"100010011101" when X = 17 AND Y = 84 else
"100010011101" when X = 18 AND Y = 84 else
"100010011101" when X = 19 AND Y = 84 else
"100010011101" when X = 20 AND Y = 84 else
"100010011101" when X = 21 AND Y = 84 else
"100010011101" when X = 22 AND Y = 84 else
"100010011101" when X = 23 AND Y = 84 else
"100010011101" when X = 24 AND Y = 84 else
"100010011101" when X = 25 AND Y = 84 else
"100010011101" when X = 26 AND Y = 84 else
"100010011101" when X = 27 AND Y = 84 else
"100010011101" when X = 28 AND Y = 84 else
"100010011101" when X = 29 AND Y = 84 else
"110111011111" when X = 30 AND Y = 84 else
"110111011111" when X = 31 AND Y = 84 else
"110111011111" when X = 32 AND Y = 84 else
"110111011111" when X = 33 AND Y = 84 else
"110111011111" when X = 34 AND Y = 84 else
"110111011111" when X = 35 AND Y = 84 else
"110111011111" when X = 36 AND Y = 84 else
"110111011111" when X = 37 AND Y = 84 else
"110111011111" when X = 38 AND Y = 84 else
"110111011111" when X = 39 AND Y = 84 else
"110111011111" when X = 40 AND Y = 84 else
"110111011111" when X = 41 AND Y = 84 else
"110111011111" when X = 42 AND Y = 84 else
"110111011111" when X = 43 AND Y = 84 else
"110111011111" when X = 44 AND Y = 84 else
"110111011111" when X = 45 AND Y = 84 else
"110111011111" when X = 46 AND Y = 84 else
"110111011111" when X = 47 AND Y = 84 else
"110111011111" when X = 48 AND Y = 84 else
"110111011111" when X = 49 AND Y = 84 else
"110111011111" when X = 50 AND Y = 84 else
"110111011111" when X = 51 AND Y = 84 else
"110111011111" when X = 52 AND Y = 84 else
"110111011111" when X = 53 AND Y = 84 else
"110111011111" when X = 54 AND Y = 84 else
"110111011111" when X = 55 AND Y = 84 else
"110111011111" when X = 56 AND Y = 84 else
"110111011111" when X = 57 AND Y = 84 else
"110111011111" when X = 58 AND Y = 84 else
"110111011111" when X = 59 AND Y = 84 else
"110111011111" when X = 60 AND Y = 84 else
"110111011111" when X = 61 AND Y = 84 else
"110111011111" when X = 62 AND Y = 84 else
"110111011111" when X = 63 AND Y = 84 else
"110111011111" when X = 64 AND Y = 84 else
"110111011111" when X = 65 AND Y = 84 else
"110111011111" when X = 66 AND Y = 84 else
"110111011111" when X = 67 AND Y = 84 else
"110111011111" when X = 68 AND Y = 84 else
"110111011111" when X = 69 AND Y = 84 else
"110111011111" when X = 70 AND Y = 84 else
"110111011111" when X = 71 AND Y = 84 else
"110111011111" when X = 72 AND Y = 84 else
"110111011111" when X = 73 AND Y = 84 else
"110111011111" when X = 74 AND Y = 84 else
"110111011111" when X = 75 AND Y = 84 else
"110111011111" when X = 76 AND Y = 84 else
"110111011111" when X = 77 AND Y = 84 else
"110111011111" when X = 78 AND Y = 84 else
"110111011111" when X = 79 AND Y = 84 else
"110111011111" when X = 80 AND Y = 84 else
"110111011111" when X = 81 AND Y = 84 else
"110111011111" when X = 82 AND Y = 84 else
"110111011111" when X = 83 AND Y = 84 else
"110111011111" when X = 84 AND Y = 84 else
"110111011111" when X = 85 AND Y = 84 else
"110111011111" when X = 86 AND Y = 84 else
"110111011111" when X = 87 AND Y = 84 else
"110111011111" when X = 88 AND Y = 84 else
"110111011111" when X = 89 AND Y = 84 else
"110111011111" when X = 90 AND Y = 84 else
"110111011111" when X = 91 AND Y = 84 else
"110111011111" when X = 92 AND Y = 84 else
"110111011111" when X = 93 AND Y = 84 else
"110111011111" when X = 94 AND Y = 84 else
"110111011111" when X = 95 AND Y = 84 else
"110111011111" when X = 96 AND Y = 84 else
"110111011111" when X = 97 AND Y = 84 else
"110111011111" when X = 98 AND Y = 84 else
"110111011111" when X = 99 AND Y = 84 else
"110111011111" when X = 100 AND Y = 84 else
"110111011111" when X = 101 AND Y = 84 else
"110111011111" when X = 102 AND Y = 84 else
"110111011111" when X = 103 AND Y = 84 else
"110111011111" when X = 104 AND Y = 84 else
"111111111111" when X = 105 AND Y = 84 else
"111111111111" when X = 106 AND Y = 84 else
"111111111111" when X = 107 AND Y = 84 else
"111111111111" when X = 108 AND Y = 84 else
"111111111111" when X = 109 AND Y = 84 else
"111111111111" when X = 110 AND Y = 84 else
"111111111111" when X = 111 AND Y = 84 else
"111111111111" when X = 112 AND Y = 84 else
"111111111111" when X = 113 AND Y = 84 else
"111111111111" when X = 114 AND Y = 84 else
"111111111111" when X = 115 AND Y = 84 else
"111111111111" when X = 116 AND Y = 84 else
"111111111111" when X = 117 AND Y = 84 else
"111111111111" when X = 118 AND Y = 84 else
"111111111111" when X = 119 AND Y = 84 else
"111111111111" when X = 120 AND Y = 84 else
"111111111111" when X = 121 AND Y = 84 else
"111111111111" when X = 122 AND Y = 84 else
"111111111111" when X = 123 AND Y = 84 else
"111111111111" when X = 124 AND Y = 84 else
"111111111111" when X = 125 AND Y = 84 else
"111111111111" when X = 126 AND Y = 84 else
"111111111111" when X = 127 AND Y = 84 else
"111111111111" when X = 128 AND Y = 84 else
"111111111111" when X = 129 AND Y = 84 else
"111111111111" when X = 130 AND Y = 84 else
"111111111111" when X = 131 AND Y = 84 else
"111111111111" when X = 132 AND Y = 84 else
"111111111111" when X = 133 AND Y = 84 else
"111111111111" when X = 134 AND Y = 84 else
"111111111111" when X = 135 AND Y = 84 else
"111111111111" when X = 136 AND Y = 84 else
"111111111111" when X = 137 AND Y = 84 else
"111111111111" when X = 138 AND Y = 84 else
"111111111111" when X = 139 AND Y = 84 else
"111111111111" when X = 140 AND Y = 84 else
"111111111111" when X = 141 AND Y = 84 else
"111111111111" when X = 142 AND Y = 84 else
"111111111111" when X = 143 AND Y = 84 else
"111111111111" when X = 144 AND Y = 84 else
"111111111111" when X = 145 AND Y = 84 else
"111111111111" when X = 146 AND Y = 84 else
"111111111111" when X = 147 AND Y = 84 else
"111111111111" when X = 148 AND Y = 84 else
"111111111111" when X = 149 AND Y = 84 else
"111111111111" when X = 150 AND Y = 84 else
"111111111111" when X = 151 AND Y = 84 else
"111111111111" when X = 152 AND Y = 84 else
"111111111111" when X = 153 AND Y = 84 else
"111111111111" when X = 154 AND Y = 84 else
"111111111111" when X = 155 AND Y = 84 else
"111111111111" when X = 156 AND Y = 84 else
"111111111111" when X = 157 AND Y = 84 else
"111111111111" when X = 158 AND Y = 84 else
"111111111111" when X = 159 AND Y = 84 else
"111111111111" when X = 160 AND Y = 84 else
"111111111111" when X = 161 AND Y = 84 else
"111111111111" when X = 162 AND Y = 84 else
"111111111111" when X = 163 AND Y = 84 else
"111111111111" when X = 164 AND Y = 84 else
"111111111111" when X = 165 AND Y = 84 else
"111111111111" when X = 166 AND Y = 84 else
"111111111111" when X = 167 AND Y = 84 else
"111111111111" when X = 168 AND Y = 84 else
"111111111111" when X = 169 AND Y = 84 else
"111111111111" when X = 170 AND Y = 84 else
"111111111111" when X = 171 AND Y = 84 else
"111111111111" when X = 172 AND Y = 84 else
"111111111111" when X = 173 AND Y = 84 else
"111111111111" when X = 174 AND Y = 84 else
"111111111111" when X = 175 AND Y = 84 else
"111111111111" when X = 176 AND Y = 84 else
"111111111111" when X = 177 AND Y = 84 else
"111111111111" when X = 178 AND Y = 84 else
"111111111111" when X = 179 AND Y = 84 else
"111111111111" when X = 180 AND Y = 84 else
"111111111111" when X = 181 AND Y = 84 else
"111111111111" when X = 182 AND Y = 84 else
"111111111111" when X = 183 AND Y = 84 else
"111111111111" when X = 184 AND Y = 84 else
"111111111111" when X = 185 AND Y = 84 else
"111111111111" when X = 186 AND Y = 84 else
"111111111111" when X = 187 AND Y = 84 else
"111111111111" when X = 188 AND Y = 84 else
"111111111111" when X = 189 AND Y = 84 else
"111111111111" when X = 190 AND Y = 84 else
"111111111111" when X = 191 AND Y = 84 else
"111111111111" when X = 192 AND Y = 84 else
"111111111111" when X = 193 AND Y = 84 else
"111111111111" when X = 194 AND Y = 84 else
"111111111111" when X = 195 AND Y = 84 else
"111111111111" when X = 196 AND Y = 84 else
"111111111111" when X = 197 AND Y = 84 else
"111111111111" when X = 198 AND Y = 84 else
"111111111111" when X = 199 AND Y = 84 else
"111111111111" when X = 200 AND Y = 84 else
"111111111111" when X = 201 AND Y = 84 else
"111111111111" when X = 202 AND Y = 84 else
"111111111111" when X = 203 AND Y = 84 else
"111111111111" when X = 204 AND Y = 84 else
"111111111111" when X = 205 AND Y = 84 else
"111111111111" when X = 206 AND Y = 84 else
"111111111111" when X = 207 AND Y = 84 else
"111111111111" when X = 208 AND Y = 84 else
"111111111111" when X = 209 AND Y = 84 else
"111111111111" when X = 210 AND Y = 84 else
"111111111111" when X = 211 AND Y = 84 else
"111111111111" when X = 212 AND Y = 84 else
"111111111111" when X = 213 AND Y = 84 else
"111111111111" when X = 214 AND Y = 84 else
"111111111111" when X = 215 AND Y = 84 else
"111111111111" when X = 216 AND Y = 84 else
"111111111111" when X = 217 AND Y = 84 else
"111111111111" when X = 218 AND Y = 84 else
"111111111111" when X = 219 AND Y = 84 else
"111111111111" when X = 220 AND Y = 84 else
"111111111111" when X = 221 AND Y = 84 else
"111111111111" when X = 222 AND Y = 84 else
"111111111111" when X = 223 AND Y = 84 else
"111111111111" when X = 224 AND Y = 84 else
"111111111111" when X = 225 AND Y = 84 else
"111111111111" when X = 226 AND Y = 84 else
"111111111111" when X = 227 AND Y = 84 else
"111111111111" when X = 228 AND Y = 84 else
"111111111111" when X = 229 AND Y = 84 else
"111111111111" when X = 230 AND Y = 84 else
"111111111111" when X = 231 AND Y = 84 else
"111111111111" when X = 232 AND Y = 84 else
"111111111111" when X = 233 AND Y = 84 else
"111111111111" when X = 234 AND Y = 84 else
"111111111111" when X = 235 AND Y = 84 else
"111111111111" when X = 236 AND Y = 84 else
"111111111111" when X = 237 AND Y = 84 else
"111111111111" when X = 238 AND Y = 84 else
"111111111111" when X = 239 AND Y = 84 else
"111111111111" when X = 240 AND Y = 84 else
"111111111111" when X = 241 AND Y = 84 else
"111111111111" when X = 242 AND Y = 84 else
"111111111111" when X = 243 AND Y = 84 else
"111111111111" when X = 244 AND Y = 84 else
"111111111111" when X = 245 AND Y = 84 else
"111111111111" when X = 246 AND Y = 84 else
"111111111111" when X = 247 AND Y = 84 else
"111111111111" when X = 248 AND Y = 84 else
"111111111111" when X = 249 AND Y = 84 else
"111111111111" when X = 250 AND Y = 84 else
"111111111111" when X = 251 AND Y = 84 else
"111111111111" when X = 252 AND Y = 84 else
"111111111111" when X = 253 AND Y = 84 else
"111111111111" when X = 254 AND Y = 84 else
"111111111111" when X = 255 AND Y = 84 else
"111111111111" when X = 256 AND Y = 84 else
"111111111111" when X = 257 AND Y = 84 else
"111111111111" when X = 258 AND Y = 84 else
"111111111111" when X = 259 AND Y = 84 else
"111111111111" when X = 260 AND Y = 84 else
"111111111111" when X = 261 AND Y = 84 else
"111111111111" when X = 262 AND Y = 84 else
"111111111111" when X = 263 AND Y = 84 else
"111111111111" when X = 264 AND Y = 84 else
"111111111111" when X = 265 AND Y = 84 else
"111111111111" when X = 266 AND Y = 84 else
"111111111111" when X = 267 AND Y = 84 else
"111111111111" when X = 268 AND Y = 84 else
"111111111111" when X = 269 AND Y = 84 else
"110111011111" when X = 270 AND Y = 84 else
"110111011111" when X = 271 AND Y = 84 else
"110111011111" when X = 272 AND Y = 84 else
"110111011111" when X = 273 AND Y = 84 else
"110111011111" when X = 274 AND Y = 84 else
"110111011111" when X = 275 AND Y = 84 else
"110111011111" when X = 276 AND Y = 84 else
"110111011111" when X = 277 AND Y = 84 else
"110111011111" when X = 278 AND Y = 84 else
"110111011111" when X = 279 AND Y = 84 else
"110111011111" when X = 280 AND Y = 84 else
"110111011111" when X = 281 AND Y = 84 else
"110111011111" when X = 282 AND Y = 84 else
"110111011111" when X = 283 AND Y = 84 else
"110111011111" when X = 284 AND Y = 84 else
"110111011111" when X = 285 AND Y = 84 else
"110111011111" when X = 286 AND Y = 84 else
"110111011111" when X = 287 AND Y = 84 else
"110111011111" when X = 288 AND Y = 84 else
"110111011111" when X = 289 AND Y = 84 else
"110111011111" when X = 290 AND Y = 84 else
"110111011111" when X = 291 AND Y = 84 else
"110111011111" when X = 292 AND Y = 84 else
"110111011111" when X = 293 AND Y = 84 else
"110111011111" when X = 294 AND Y = 84 else
"110111011111" when X = 295 AND Y = 84 else
"110111011111" when X = 296 AND Y = 84 else
"110111011111" when X = 297 AND Y = 84 else
"110111011111" when X = 298 AND Y = 84 else
"110111011111" when X = 299 AND Y = 84 else
"110111011111" when X = 300 AND Y = 84 else
"110111011111" when X = 301 AND Y = 84 else
"110111011111" when X = 302 AND Y = 84 else
"110111011111" when X = 303 AND Y = 84 else
"110111011111" when X = 304 AND Y = 84 else
"110111011111" when X = 305 AND Y = 84 else
"110111011111" when X = 306 AND Y = 84 else
"110111011111" when X = 307 AND Y = 84 else
"110111011111" when X = 308 AND Y = 84 else
"110111011111" when X = 309 AND Y = 84 else
"110111011111" when X = 310 AND Y = 84 else
"110111011111" when X = 311 AND Y = 84 else
"110111011111" when X = 312 AND Y = 84 else
"110111011111" when X = 313 AND Y = 84 else
"110111011111" when X = 314 AND Y = 84 else
"110111011111" when X = 315 AND Y = 84 else
"110111011111" when X = 316 AND Y = 84 else
"110111011111" when X = 317 AND Y = 84 else
"110111011111" when X = 318 AND Y = 84 else
"110111011111" when X = 319 AND Y = 84 else
"000000000000" when X = 320 AND Y = 84 else
"000000000000" when X = 321 AND Y = 84 else
"000000000000" when X = 322 AND Y = 84 else
"000000000000" when X = 323 AND Y = 84 else
"000000000000" when X = 324 AND Y = 84 else
"100010011101" when X = 0 AND Y = 85 else
"100010011101" when X = 1 AND Y = 85 else
"100010011101" when X = 2 AND Y = 85 else
"100010011101" when X = 3 AND Y = 85 else
"100010011101" when X = 4 AND Y = 85 else
"100010011101" when X = 5 AND Y = 85 else
"100010011101" when X = 6 AND Y = 85 else
"100010011101" when X = 7 AND Y = 85 else
"100010011101" when X = 8 AND Y = 85 else
"100010011101" when X = 9 AND Y = 85 else
"100010011101" when X = 10 AND Y = 85 else
"100010011101" when X = 11 AND Y = 85 else
"100010011101" when X = 12 AND Y = 85 else
"100010011101" when X = 13 AND Y = 85 else
"100010011101" when X = 14 AND Y = 85 else
"100010011101" when X = 15 AND Y = 85 else
"100010011101" when X = 16 AND Y = 85 else
"100010011101" when X = 17 AND Y = 85 else
"100010011101" when X = 18 AND Y = 85 else
"100010011101" when X = 19 AND Y = 85 else
"100010011101" when X = 20 AND Y = 85 else
"100010011101" when X = 21 AND Y = 85 else
"100010011101" when X = 22 AND Y = 85 else
"100010011101" when X = 23 AND Y = 85 else
"100010011101" when X = 24 AND Y = 85 else
"110111011111" when X = 25 AND Y = 85 else
"110111011111" when X = 26 AND Y = 85 else
"110111011111" when X = 27 AND Y = 85 else
"110111011111" when X = 28 AND Y = 85 else
"110111011111" when X = 29 AND Y = 85 else
"110111011111" when X = 30 AND Y = 85 else
"110111011111" when X = 31 AND Y = 85 else
"110111011111" when X = 32 AND Y = 85 else
"110111011111" when X = 33 AND Y = 85 else
"110111011111" when X = 34 AND Y = 85 else
"110111011111" when X = 35 AND Y = 85 else
"110111011111" when X = 36 AND Y = 85 else
"110111011111" when X = 37 AND Y = 85 else
"110111011111" when X = 38 AND Y = 85 else
"110111011111" when X = 39 AND Y = 85 else
"110111011111" when X = 40 AND Y = 85 else
"110111011111" when X = 41 AND Y = 85 else
"110111011111" when X = 42 AND Y = 85 else
"110111011111" when X = 43 AND Y = 85 else
"110111011111" when X = 44 AND Y = 85 else
"110111011111" when X = 45 AND Y = 85 else
"110111011111" when X = 46 AND Y = 85 else
"110111011111" when X = 47 AND Y = 85 else
"110111011111" when X = 48 AND Y = 85 else
"110111011111" when X = 49 AND Y = 85 else
"110111011111" when X = 50 AND Y = 85 else
"110111011111" when X = 51 AND Y = 85 else
"110111011111" when X = 52 AND Y = 85 else
"110111011111" when X = 53 AND Y = 85 else
"110111011111" when X = 54 AND Y = 85 else
"110111011111" when X = 55 AND Y = 85 else
"110111011111" when X = 56 AND Y = 85 else
"110111011111" when X = 57 AND Y = 85 else
"110111011111" when X = 58 AND Y = 85 else
"110111011111" when X = 59 AND Y = 85 else
"110111011111" when X = 60 AND Y = 85 else
"110111011111" when X = 61 AND Y = 85 else
"110111011111" when X = 62 AND Y = 85 else
"110111011111" when X = 63 AND Y = 85 else
"110111011111" when X = 64 AND Y = 85 else
"110111011111" when X = 65 AND Y = 85 else
"110111011111" when X = 66 AND Y = 85 else
"110111011111" when X = 67 AND Y = 85 else
"110111011111" when X = 68 AND Y = 85 else
"110111011111" when X = 69 AND Y = 85 else
"110111011111" when X = 70 AND Y = 85 else
"110111011111" when X = 71 AND Y = 85 else
"110111011111" when X = 72 AND Y = 85 else
"110111011111" when X = 73 AND Y = 85 else
"110111011111" when X = 74 AND Y = 85 else
"110111011111" when X = 75 AND Y = 85 else
"110111011111" when X = 76 AND Y = 85 else
"110111011111" when X = 77 AND Y = 85 else
"110111011111" when X = 78 AND Y = 85 else
"110111011111" when X = 79 AND Y = 85 else
"110111011111" when X = 80 AND Y = 85 else
"110111011111" when X = 81 AND Y = 85 else
"110111011111" when X = 82 AND Y = 85 else
"110111011111" when X = 83 AND Y = 85 else
"110111011111" when X = 84 AND Y = 85 else
"110111011111" when X = 85 AND Y = 85 else
"110111011111" when X = 86 AND Y = 85 else
"110111011111" when X = 87 AND Y = 85 else
"110111011111" when X = 88 AND Y = 85 else
"110111011111" when X = 89 AND Y = 85 else
"110111011111" when X = 90 AND Y = 85 else
"110111011111" when X = 91 AND Y = 85 else
"110111011111" when X = 92 AND Y = 85 else
"110111011111" when X = 93 AND Y = 85 else
"110111011111" when X = 94 AND Y = 85 else
"110111011111" when X = 95 AND Y = 85 else
"110111011111" when X = 96 AND Y = 85 else
"110111011111" when X = 97 AND Y = 85 else
"110111011111" when X = 98 AND Y = 85 else
"110111011111" when X = 99 AND Y = 85 else
"111111111111" when X = 100 AND Y = 85 else
"111111111111" when X = 101 AND Y = 85 else
"111111111111" when X = 102 AND Y = 85 else
"111111111111" when X = 103 AND Y = 85 else
"111111111111" when X = 104 AND Y = 85 else
"111111111111" when X = 105 AND Y = 85 else
"111111111111" when X = 106 AND Y = 85 else
"111111111111" when X = 107 AND Y = 85 else
"111111111111" when X = 108 AND Y = 85 else
"111111111111" when X = 109 AND Y = 85 else
"111111111111" when X = 110 AND Y = 85 else
"111111111111" when X = 111 AND Y = 85 else
"111111111111" when X = 112 AND Y = 85 else
"111111111111" when X = 113 AND Y = 85 else
"111111111111" when X = 114 AND Y = 85 else
"111111111111" when X = 115 AND Y = 85 else
"111111111111" when X = 116 AND Y = 85 else
"111111111111" when X = 117 AND Y = 85 else
"111111111111" when X = 118 AND Y = 85 else
"111111111111" when X = 119 AND Y = 85 else
"111111111111" when X = 120 AND Y = 85 else
"111111111111" when X = 121 AND Y = 85 else
"111111111111" when X = 122 AND Y = 85 else
"111111111111" when X = 123 AND Y = 85 else
"111111111111" when X = 124 AND Y = 85 else
"111111111111" when X = 125 AND Y = 85 else
"111111111111" when X = 126 AND Y = 85 else
"111111111111" when X = 127 AND Y = 85 else
"111111111111" when X = 128 AND Y = 85 else
"111111111111" when X = 129 AND Y = 85 else
"111111111111" when X = 130 AND Y = 85 else
"111111111111" when X = 131 AND Y = 85 else
"111111111111" when X = 132 AND Y = 85 else
"111111111111" when X = 133 AND Y = 85 else
"111111111111" when X = 134 AND Y = 85 else
"111111111111" when X = 135 AND Y = 85 else
"111111111111" when X = 136 AND Y = 85 else
"111111111111" when X = 137 AND Y = 85 else
"111111111111" when X = 138 AND Y = 85 else
"111111111111" when X = 139 AND Y = 85 else
"111111111111" when X = 140 AND Y = 85 else
"111111111111" when X = 141 AND Y = 85 else
"111111111111" when X = 142 AND Y = 85 else
"111111111111" when X = 143 AND Y = 85 else
"111111111111" when X = 144 AND Y = 85 else
"111111111111" when X = 145 AND Y = 85 else
"111111111111" when X = 146 AND Y = 85 else
"111111111111" when X = 147 AND Y = 85 else
"111111111111" when X = 148 AND Y = 85 else
"111111111111" when X = 149 AND Y = 85 else
"111111111111" when X = 150 AND Y = 85 else
"111111111111" when X = 151 AND Y = 85 else
"111111111111" when X = 152 AND Y = 85 else
"111111111111" when X = 153 AND Y = 85 else
"111111111111" when X = 154 AND Y = 85 else
"111111111111" when X = 155 AND Y = 85 else
"111111111111" when X = 156 AND Y = 85 else
"111111111111" when X = 157 AND Y = 85 else
"111111111111" when X = 158 AND Y = 85 else
"111111111111" when X = 159 AND Y = 85 else
"111111111111" when X = 160 AND Y = 85 else
"111111111111" when X = 161 AND Y = 85 else
"111111111111" when X = 162 AND Y = 85 else
"111111111111" when X = 163 AND Y = 85 else
"111111111111" when X = 164 AND Y = 85 else
"111111111111" when X = 165 AND Y = 85 else
"111111111111" when X = 166 AND Y = 85 else
"111111111111" when X = 167 AND Y = 85 else
"111111111111" when X = 168 AND Y = 85 else
"111111111111" when X = 169 AND Y = 85 else
"111111111111" when X = 170 AND Y = 85 else
"111111111111" when X = 171 AND Y = 85 else
"111111111111" when X = 172 AND Y = 85 else
"111111111111" when X = 173 AND Y = 85 else
"111111111111" when X = 174 AND Y = 85 else
"111111111111" when X = 175 AND Y = 85 else
"111111111111" when X = 176 AND Y = 85 else
"111111111111" when X = 177 AND Y = 85 else
"111111111111" when X = 178 AND Y = 85 else
"111111111111" when X = 179 AND Y = 85 else
"111111111111" when X = 180 AND Y = 85 else
"111111111111" when X = 181 AND Y = 85 else
"111111111111" when X = 182 AND Y = 85 else
"111111111111" when X = 183 AND Y = 85 else
"111111111111" when X = 184 AND Y = 85 else
"111111111111" when X = 185 AND Y = 85 else
"111111111111" when X = 186 AND Y = 85 else
"111111111111" when X = 187 AND Y = 85 else
"111111111111" when X = 188 AND Y = 85 else
"111111111111" when X = 189 AND Y = 85 else
"111111111111" when X = 190 AND Y = 85 else
"111111111111" when X = 191 AND Y = 85 else
"111111111111" when X = 192 AND Y = 85 else
"111111111111" when X = 193 AND Y = 85 else
"111111111111" when X = 194 AND Y = 85 else
"111111111111" when X = 195 AND Y = 85 else
"111111111111" when X = 196 AND Y = 85 else
"111111111111" when X = 197 AND Y = 85 else
"111111111111" when X = 198 AND Y = 85 else
"111111111111" when X = 199 AND Y = 85 else
"111111111111" when X = 200 AND Y = 85 else
"111111111111" when X = 201 AND Y = 85 else
"111111111111" when X = 202 AND Y = 85 else
"111111111111" when X = 203 AND Y = 85 else
"111111111111" when X = 204 AND Y = 85 else
"111111111111" when X = 205 AND Y = 85 else
"111111111111" when X = 206 AND Y = 85 else
"111111111111" when X = 207 AND Y = 85 else
"111111111111" when X = 208 AND Y = 85 else
"111111111111" when X = 209 AND Y = 85 else
"111111111111" when X = 210 AND Y = 85 else
"111111111111" when X = 211 AND Y = 85 else
"111111111111" when X = 212 AND Y = 85 else
"111111111111" when X = 213 AND Y = 85 else
"111111111111" when X = 214 AND Y = 85 else
"111111111111" when X = 215 AND Y = 85 else
"111111111111" when X = 216 AND Y = 85 else
"111111111111" when X = 217 AND Y = 85 else
"111111111111" when X = 218 AND Y = 85 else
"111111111111" when X = 219 AND Y = 85 else
"111111111111" when X = 220 AND Y = 85 else
"111111111111" when X = 221 AND Y = 85 else
"111111111111" when X = 222 AND Y = 85 else
"111111111111" when X = 223 AND Y = 85 else
"111111111111" when X = 224 AND Y = 85 else
"111111111111" when X = 225 AND Y = 85 else
"111111111111" when X = 226 AND Y = 85 else
"111111111111" when X = 227 AND Y = 85 else
"111111111111" when X = 228 AND Y = 85 else
"111111111111" when X = 229 AND Y = 85 else
"111111111111" when X = 230 AND Y = 85 else
"111111111111" when X = 231 AND Y = 85 else
"111111111111" when X = 232 AND Y = 85 else
"111111111111" when X = 233 AND Y = 85 else
"111111111111" when X = 234 AND Y = 85 else
"111111111111" when X = 235 AND Y = 85 else
"111111111111" when X = 236 AND Y = 85 else
"111111111111" when X = 237 AND Y = 85 else
"111111111111" when X = 238 AND Y = 85 else
"111111111111" when X = 239 AND Y = 85 else
"111111111111" when X = 240 AND Y = 85 else
"111111111111" when X = 241 AND Y = 85 else
"111111111111" when X = 242 AND Y = 85 else
"111111111111" when X = 243 AND Y = 85 else
"111111111111" when X = 244 AND Y = 85 else
"111111111111" when X = 245 AND Y = 85 else
"111111111111" when X = 246 AND Y = 85 else
"111111111111" when X = 247 AND Y = 85 else
"111111111111" when X = 248 AND Y = 85 else
"111111111111" when X = 249 AND Y = 85 else
"111111111111" when X = 250 AND Y = 85 else
"111111111111" when X = 251 AND Y = 85 else
"111111111111" when X = 252 AND Y = 85 else
"111111111111" when X = 253 AND Y = 85 else
"111111111111" when X = 254 AND Y = 85 else
"111111111111" when X = 255 AND Y = 85 else
"111111111111" when X = 256 AND Y = 85 else
"111111111111" when X = 257 AND Y = 85 else
"111111111111" when X = 258 AND Y = 85 else
"111111111111" when X = 259 AND Y = 85 else
"111111111111" when X = 260 AND Y = 85 else
"111111111111" when X = 261 AND Y = 85 else
"111111111111" when X = 262 AND Y = 85 else
"111111111111" when X = 263 AND Y = 85 else
"111111111111" when X = 264 AND Y = 85 else
"111111111111" when X = 265 AND Y = 85 else
"111111111111" when X = 266 AND Y = 85 else
"111111111111" when X = 267 AND Y = 85 else
"111111111111" when X = 268 AND Y = 85 else
"111111111111" when X = 269 AND Y = 85 else
"111111111111" when X = 270 AND Y = 85 else
"111111111111" when X = 271 AND Y = 85 else
"111111111111" when X = 272 AND Y = 85 else
"111111111111" when X = 273 AND Y = 85 else
"111111111111" when X = 274 AND Y = 85 else
"110111011111" when X = 275 AND Y = 85 else
"110111011111" when X = 276 AND Y = 85 else
"110111011111" when X = 277 AND Y = 85 else
"110111011111" when X = 278 AND Y = 85 else
"110111011111" when X = 279 AND Y = 85 else
"110111011111" when X = 280 AND Y = 85 else
"110111011111" when X = 281 AND Y = 85 else
"110111011111" when X = 282 AND Y = 85 else
"110111011111" when X = 283 AND Y = 85 else
"110111011111" when X = 284 AND Y = 85 else
"110111011111" when X = 285 AND Y = 85 else
"110111011111" when X = 286 AND Y = 85 else
"110111011111" when X = 287 AND Y = 85 else
"110111011111" when X = 288 AND Y = 85 else
"110111011111" when X = 289 AND Y = 85 else
"110111011111" when X = 290 AND Y = 85 else
"110111011111" when X = 291 AND Y = 85 else
"110111011111" when X = 292 AND Y = 85 else
"110111011111" when X = 293 AND Y = 85 else
"110111011111" when X = 294 AND Y = 85 else
"110111011111" when X = 295 AND Y = 85 else
"110111011111" when X = 296 AND Y = 85 else
"110111011111" when X = 297 AND Y = 85 else
"110111011111" when X = 298 AND Y = 85 else
"110111011111" when X = 299 AND Y = 85 else
"110111011111" when X = 300 AND Y = 85 else
"110111011111" when X = 301 AND Y = 85 else
"110111011111" when X = 302 AND Y = 85 else
"110111011111" when X = 303 AND Y = 85 else
"110111011111" when X = 304 AND Y = 85 else
"110111011111" when X = 305 AND Y = 85 else
"110111011111" when X = 306 AND Y = 85 else
"110111011111" when X = 307 AND Y = 85 else
"110111011111" when X = 308 AND Y = 85 else
"110111011111" when X = 309 AND Y = 85 else
"110111011111" when X = 310 AND Y = 85 else
"110111011111" when X = 311 AND Y = 85 else
"110111011111" when X = 312 AND Y = 85 else
"110111011111" when X = 313 AND Y = 85 else
"110111011111" when X = 314 AND Y = 85 else
"110111011111" when X = 315 AND Y = 85 else
"110111011111" when X = 316 AND Y = 85 else
"110111011111" when X = 317 AND Y = 85 else
"110111011111" when X = 318 AND Y = 85 else
"110111011111" when X = 319 AND Y = 85 else
"000000000000" when X = 320 AND Y = 85 else
"000000000000" when X = 321 AND Y = 85 else
"000000000000" when X = 322 AND Y = 85 else
"000000000000" when X = 323 AND Y = 85 else
"000000000000" when X = 324 AND Y = 85 else
"100010011101" when X = 0 AND Y = 86 else
"100010011101" when X = 1 AND Y = 86 else
"100010011101" when X = 2 AND Y = 86 else
"100010011101" when X = 3 AND Y = 86 else
"100010011101" when X = 4 AND Y = 86 else
"100010011101" when X = 5 AND Y = 86 else
"100010011101" when X = 6 AND Y = 86 else
"100010011101" when X = 7 AND Y = 86 else
"100010011101" when X = 8 AND Y = 86 else
"100010011101" when X = 9 AND Y = 86 else
"100010011101" when X = 10 AND Y = 86 else
"100010011101" when X = 11 AND Y = 86 else
"100010011101" when X = 12 AND Y = 86 else
"100010011101" when X = 13 AND Y = 86 else
"100010011101" when X = 14 AND Y = 86 else
"100010011101" when X = 15 AND Y = 86 else
"100010011101" when X = 16 AND Y = 86 else
"100010011101" when X = 17 AND Y = 86 else
"100010011101" when X = 18 AND Y = 86 else
"100010011101" when X = 19 AND Y = 86 else
"100010011101" when X = 20 AND Y = 86 else
"100010011101" when X = 21 AND Y = 86 else
"100010011101" when X = 22 AND Y = 86 else
"100010011101" when X = 23 AND Y = 86 else
"100010011101" when X = 24 AND Y = 86 else
"110111011111" when X = 25 AND Y = 86 else
"110111011111" when X = 26 AND Y = 86 else
"110111011111" when X = 27 AND Y = 86 else
"110111011111" when X = 28 AND Y = 86 else
"110111011111" when X = 29 AND Y = 86 else
"110111011111" when X = 30 AND Y = 86 else
"110111011111" when X = 31 AND Y = 86 else
"110111011111" when X = 32 AND Y = 86 else
"110111011111" when X = 33 AND Y = 86 else
"110111011111" when X = 34 AND Y = 86 else
"110111011111" when X = 35 AND Y = 86 else
"110111011111" when X = 36 AND Y = 86 else
"110111011111" when X = 37 AND Y = 86 else
"110111011111" when X = 38 AND Y = 86 else
"110111011111" when X = 39 AND Y = 86 else
"110111011111" when X = 40 AND Y = 86 else
"110111011111" when X = 41 AND Y = 86 else
"110111011111" when X = 42 AND Y = 86 else
"110111011111" when X = 43 AND Y = 86 else
"110111011111" when X = 44 AND Y = 86 else
"110111011111" when X = 45 AND Y = 86 else
"110111011111" when X = 46 AND Y = 86 else
"110111011111" when X = 47 AND Y = 86 else
"110111011111" when X = 48 AND Y = 86 else
"110111011111" when X = 49 AND Y = 86 else
"110111011111" when X = 50 AND Y = 86 else
"110111011111" when X = 51 AND Y = 86 else
"110111011111" when X = 52 AND Y = 86 else
"110111011111" when X = 53 AND Y = 86 else
"110111011111" when X = 54 AND Y = 86 else
"110111011111" when X = 55 AND Y = 86 else
"110111011111" when X = 56 AND Y = 86 else
"110111011111" when X = 57 AND Y = 86 else
"110111011111" when X = 58 AND Y = 86 else
"110111011111" when X = 59 AND Y = 86 else
"110111011111" when X = 60 AND Y = 86 else
"110111011111" when X = 61 AND Y = 86 else
"110111011111" when X = 62 AND Y = 86 else
"110111011111" when X = 63 AND Y = 86 else
"110111011111" when X = 64 AND Y = 86 else
"110111011111" when X = 65 AND Y = 86 else
"110111011111" when X = 66 AND Y = 86 else
"110111011111" when X = 67 AND Y = 86 else
"110111011111" when X = 68 AND Y = 86 else
"110111011111" when X = 69 AND Y = 86 else
"110111011111" when X = 70 AND Y = 86 else
"110111011111" when X = 71 AND Y = 86 else
"110111011111" when X = 72 AND Y = 86 else
"110111011111" when X = 73 AND Y = 86 else
"110111011111" when X = 74 AND Y = 86 else
"110111011111" when X = 75 AND Y = 86 else
"110111011111" when X = 76 AND Y = 86 else
"110111011111" when X = 77 AND Y = 86 else
"110111011111" when X = 78 AND Y = 86 else
"110111011111" when X = 79 AND Y = 86 else
"110111011111" when X = 80 AND Y = 86 else
"110111011111" when X = 81 AND Y = 86 else
"110111011111" when X = 82 AND Y = 86 else
"110111011111" when X = 83 AND Y = 86 else
"110111011111" when X = 84 AND Y = 86 else
"110111011111" when X = 85 AND Y = 86 else
"110111011111" when X = 86 AND Y = 86 else
"110111011111" when X = 87 AND Y = 86 else
"110111011111" when X = 88 AND Y = 86 else
"110111011111" when X = 89 AND Y = 86 else
"110111011111" when X = 90 AND Y = 86 else
"110111011111" when X = 91 AND Y = 86 else
"110111011111" when X = 92 AND Y = 86 else
"110111011111" when X = 93 AND Y = 86 else
"110111011111" when X = 94 AND Y = 86 else
"110111011111" when X = 95 AND Y = 86 else
"110111011111" when X = 96 AND Y = 86 else
"110111011111" when X = 97 AND Y = 86 else
"110111011111" when X = 98 AND Y = 86 else
"110111011111" when X = 99 AND Y = 86 else
"111111111111" when X = 100 AND Y = 86 else
"111111111111" when X = 101 AND Y = 86 else
"111111111111" when X = 102 AND Y = 86 else
"111111111111" when X = 103 AND Y = 86 else
"111111111111" when X = 104 AND Y = 86 else
"111111111111" when X = 105 AND Y = 86 else
"111111111111" when X = 106 AND Y = 86 else
"111111111111" when X = 107 AND Y = 86 else
"111111111111" when X = 108 AND Y = 86 else
"111111111111" when X = 109 AND Y = 86 else
"111111111111" when X = 110 AND Y = 86 else
"111111111111" when X = 111 AND Y = 86 else
"111111111111" when X = 112 AND Y = 86 else
"111111111111" when X = 113 AND Y = 86 else
"111111111111" when X = 114 AND Y = 86 else
"111111111111" when X = 115 AND Y = 86 else
"111111111111" when X = 116 AND Y = 86 else
"111111111111" when X = 117 AND Y = 86 else
"111111111111" when X = 118 AND Y = 86 else
"111111111111" when X = 119 AND Y = 86 else
"111111111111" when X = 120 AND Y = 86 else
"111111111111" when X = 121 AND Y = 86 else
"111111111111" when X = 122 AND Y = 86 else
"111111111111" when X = 123 AND Y = 86 else
"111111111111" when X = 124 AND Y = 86 else
"111111111111" when X = 125 AND Y = 86 else
"111111111111" when X = 126 AND Y = 86 else
"111111111111" when X = 127 AND Y = 86 else
"111111111111" when X = 128 AND Y = 86 else
"111111111111" when X = 129 AND Y = 86 else
"111111111111" when X = 130 AND Y = 86 else
"111111111111" when X = 131 AND Y = 86 else
"111111111111" when X = 132 AND Y = 86 else
"111111111111" when X = 133 AND Y = 86 else
"111111111111" when X = 134 AND Y = 86 else
"111111111111" when X = 135 AND Y = 86 else
"111111111111" when X = 136 AND Y = 86 else
"111111111111" when X = 137 AND Y = 86 else
"111111111111" when X = 138 AND Y = 86 else
"111111111111" when X = 139 AND Y = 86 else
"111111111111" when X = 140 AND Y = 86 else
"111111111111" when X = 141 AND Y = 86 else
"111111111111" when X = 142 AND Y = 86 else
"111111111111" when X = 143 AND Y = 86 else
"111111111111" when X = 144 AND Y = 86 else
"111111111111" when X = 145 AND Y = 86 else
"111111111111" when X = 146 AND Y = 86 else
"111111111111" when X = 147 AND Y = 86 else
"111111111111" when X = 148 AND Y = 86 else
"111111111111" when X = 149 AND Y = 86 else
"111111111111" when X = 150 AND Y = 86 else
"111111111111" when X = 151 AND Y = 86 else
"111111111111" when X = 152 AND Y = 86 else
"111111111111" when X = 153 AND Y = 86 else
"111111111111" when X = 154 AND Y = 86 else
"111111111111" when X = 155 AND Y = 86 else
"111111111111" when X = 156 AND Y = 86 else
"111111111111" when X = 157 AND Y = 86 else
"111111111111" when X = 158 AND Y = 86 else
"111111111111" when X = 159 AND Y = 86 else
"111111111111" when X = 160 AND Y = 86 else
"111111111111" when X = 161 AND Y = 86 else
"111111111111" when X = 162 AND Y = 86 else
"111111111111" when X = 163 AND Y = 86 else
"111111111111" when X = 164 AND Y = 86 else
"111111111111" when X = 165 AND Y = 86 else
"111111111111" when X = 166 AND Y = 86 else
"111111111111" when X = 167 AND Y = 86 else
"111111111111" when X = 168 AND Y = 86 else
"111111111111" when X = 169 AND Y = 86 else
"111111111111" when X = 170 AND Y = 86 else
"111111111111" when X = 171 AND Y = 86 else
"111111111111" when X = 172 AND Y = 86 else
"111111111111" when X = 173 AND Y = 86 else
"111111111111" when X = 174 AND Y = 86 else
"111111111111" when X = 175 AND Y = 86 else
"111111111111" when X = 176 AND Y = 86 else
"111111111111" when X = 177 AND Y = 86 else
"111111111111" when X = 178 AND Y = 86 else
"111111111111" when X = 179 AND Y = 86 else
"111111111111" when X = 180 AND Y = 86 else
"111111111111" when X = 181 AND Y = 86 else
"111111111111" when X = 182 AND Y = 86 else
"111111111111" when X = 183 AND Y = 86 else
"111111111111" when X = 184 AND Y = 86 else
"111111111111" when X = 185 AND Y = 86 else
"111111111111" when X = 186 AND Y = 86 else
"111111111111" when X = 187 AND Y = 86 else
"111111111111" when X = 188 AND Y = 86 else
"111111111111" when X = 189 AND Y = 86 else
"111111111111" when X = 190 AND Y = 86 else
"111111111111" when X = 191 AND Y = 86 else
"111111111111" when X = 192 AND Y = 86 else
"111111111111" when X = 193 AND Y = 86 else
"111111111111" when X = 194 AND Y = 86 else
"111111111111" when X = 195 AND Y = 86 else
"111111111111" when X = 196 AND Y = 86 else
"111111111111" when X = 197 AND Y = 86 else
"111111111111" when X = 198 AND Y = 86 else
"111111111111" when X = 199 AND Y = 86 else
"111111111111" when X = 200 AND Y = 86 else
"111111111111" when X = 201 AND Y = 86 else
"111111111111" when X = 202 AND Y = 86 else
"111111111111" when X = 203 AND Y = 86 else
"111111111111" when X = 204 AND Y = 86 else
"111111111111" when X = 205 AND Y = 86 else
"111111111111" when X = 206 AND Y = 86 else
"111111111111" when X = 207 AND Y = 86 else
"111111111111" when X = 208 AND Y = 86 else
"111111111111" when X = 209 AND Y = 86 else
"111111111111" when X = 210 AND Y = 86 else
"111111111111" when X = 211 AND Y = 86 else
"111111111111" when X = 212 AND Y = 86 else
"111111111111" when X = 213 AND Y = 86 else
"111111111111" when X = 214 AND Y = 86 else
"111111111111" when X = 215 AND Y = 86 else
"111111111111" when X = 216 AND Y = 86 else
"111111111111" when X = 217 AND Y = 86 else
"111111111111" when X = 218 AND Y = 86 else
"111111111111" when X = 219 AND Y = 86 else
"111111111111" when X = 220 AND Y = 86 else
"111111111111" when X = 221 AND Y = 86 else
"111111111111" when X = 222 AND Y = 86 else
"111111111111" when X = 223 AND Y = 86 else
"111111111111" when X = 224 AND Y = 86 else
"111111111111" when X = 225 AND Y = 86 else
"111111111111" when X = 226 AND Y = 86 else
"111111111111" when X = 227 AND Y = 86 else
"111111111111" when X = 228 AND Y = 86 else
"111111111111" when X = 229 AND Y = 86 else
"111111111111" when X = 230 AND Y = 86 else
"111111111111" when X = 231 AND Y = 86 else
"111111111111" when X = 232 AND Y = 86 else
"111111111111" when X = 233 AND Y = 86 else
"111111111111" when X = 234 AND Y = 86 else
"111111111111" when X = 235 AND Y = 86 else
"111111111111" when X = 236 AND Y = 86 else
"111111111111" when X = 237 AND Y = 86 else
"111111111111" when X = 238 AND Y = 86 else
"111111111111" when X = 239 AND Y = 86 else
"111111111111" when X = 240 AND Y = 86 else
"111111111111" when X = 241 AND Y = 86 else
"111111111111" when X = 242 AND Y = 86 else
"111111111111" when X = 243 AND Y = 86 else
"111111111111" when X = 244 AND Y = 86 else
"111111111111" when X = 245 AND Y = 86 else
"111111111111" when X = 246 AND Y = 86 else
"111111111111" when X = 247 AND Y = 86 else
"111111111111" when X = 248 AND Y = 86 else
"111111111111" when X = 249 AND Y = 86 else
"111111111111" when X = 250 AND Y = 86 else
"111111111111" when X = 251 AND Y = 86 else
"111111111111" when X = 252 AND Y = 86 else
"111111111111" when X = 253 AND Y = 86 else
"111111111111" when X = 254 AND Y = 86 else
"111111111111" when X = 255 AND Y = 86 else
"111111111111" when X = 256 AND Y = 86 else
"111111111111" when X = 257 AND Y = 86 else
"111111111111" when X = 258 AND Y = 86 else
"111111111111" when X = 259 AND Y = 86 else
"111111111111" when X = 260 AND Y = 86 else
"111111111111" when X = 261 AND Y = 86 else
"111111111111" when X = 262 AND Y = 86 else
"111111111111" when X = 263 AND Y = 86 else
"111111111111" when X = 264 AND Y = 86 else
"111111111111" when X = 265 AND Y = 86 else
"111111111111" when X = 266 AND Y = 86 else
"111111111111" when X = 267 AND Y = 86 else
"111111111111" when X = 268 AND Y = 86 else
"111111111111" when X = 269 AND Y = 86 else
"111111111111" when X = 270 AND Y = 86 else
"111111111111" when X = 271 AND Y = 86 else
"111111111111" when X = 272 AND Y = 86 else
"111111111111" when X = 273 AND Y = 86 else
"111111111111" when X = 274 AND Y = 86 else
"110111011111" when X = 275 AND Y = 86 else
"110111011111" when X = 276 AND Y = 86 else
"110111011111" when X = 277 AND Y = 86 else
"110111011111" when X = 278 AND Y = 86 else
"110111011111" when X = 279 AND Y = 86 else
"110111011111" when X = 280 AND Y = 86 else
"110111011111" when X = 281 AND Y = 86 else
"110111011111" when X = 282 AND Y = 86 else
"110111011111" when X = 283 AND Y = 86 else
"110111011111" when X = 284 AND Y = 86 else
"110111011111" when X = 285 AND Y = 86 else
"110111011111" when X = 286 AND Y = 86 else
"110111011111" when X = 287 AND Y = 86 else
"110111011111" when X = 288 AND Y = 86 else
"110111011111" when X = 289 AND Y = 86 else
"110111011111" when X = 290 AND Y = 86 else
"110111011111" when X = 291 AND Y = 86 else
"110111011111" when X = 292 AND Y = 86 else
"110111011111" when X = 293 AND Y = 86 else
"110111011111" when X = 294 AND Y = 86 else
"110111011111" when X = 295 AND Y = 86 else
"110111011111" when X = 296 AND Y = 86 else
"110111011111" when X = 297 AND Y = 86 else
"110111011111" when X = 298 AND Y = 86 else
"110111011111" when X = 299 AND Y = 86 else
"110111011111" when X = 300 AND Y = 86 else
"110111011111" when X = 301 AND Y = 86 else
"110111011111" when X = 302 AND Y = 86 else
"110111011111" when X = 303 AND Y = 86 else
"110111011111" when X = 304 AND Y = 86 else
"110111011111" when X = 305 AND Y = 86 else
"110111011111" when X = 306 AND Y = 86 else
"110111011111" when X = 307 AND Y = 86 else
"110111011111" when X = 308 AND Y = 86 else
"110111011111" when X = 309 AND Y = 86 else
"110111011111" when X = 310 AND Y = 86 else
"110111011111" when X = 311 AND Y = 86 else
"110111011111" when X = 312 AND Y = 86 else
"110111011111" when X = 313 AND Y = 86 else
"110111011111" when X = 314 AND Y = 86 else
"110111011111" when X = 315 AND Y = 86 else
"110111011111" when X = 316 AND Y = 86 else
"110111011111" when X = 317 AND Y = 86 else
"110111011111" when X = 318 AND Y = 86 else
"110111011111" when X = 319 AND Y = 86 else
"000000000000" when X = 320 AND Y = 86 else
"000000000000" when X = 321 AND Y = 86 else
"000000000000" when X = 322 AND Y = 86 else
"000000000000" when X = 323 AND Y = 86 else
"000000000000" when X = 324 AND Y = 86 else
"100010011101" when X = 0 AND Y = 87 else
"100010011101" when X = 1 AND Y = 87 else
"100010011101" when X = 2 AND Y = 87 else
"100010011101" when X = 3 AND Y = 87 else
"100010011101" when X = 4 AND Y = 87 else
"100010011101" when X = 5 AND Y = 87 else
"100010011101" when X = 6 AND Y = 87 else
"100010011101" when X = 7 AND Y = 87 else
"100010011101" when X = 8 AND Y = 87 else
"100010011101" when X = 9 AND Y = 87 else
"100010011101" when X = 10 AND Y = 87 else
"100010011101" when X = 11 AND Y = 87 else
"100010011101" when X = 12 AND Y = 87 else
"100010011101" when X = 13 AND Y = 87 else
"100010011101" when X = 14 AND Y = 87 else
"100010011101" when X = 15 AND Y = 87 else
"100010011101" when X = 16 AND Y = 87 else
"100010011101" when X = 17 AND Y = 87 else
"100010011101" when X = 18 AND Y = 87 else
"100010011101" when X = 19 AND Y = 87 else
"100010011101" when X = 20 AND Y = 87 else
"100010011101" when X = 21 AND Y = 87 else
"100010011101" when X = 22 AND Y = 87 else
"100010011101" when X = 23 AND Y = 87 else
"100010011101" when X = 24 AND Y = 87 else
"110111011111" when X = 25 AND Y = 87 else
"110111011111" when X = 26 AND Y = 87 else
"110111011111" when X = 27 AND Y = 87 else
"110111011111" when X = 28 AND Y = 87 else
"110111011111" when X = 29 AND Y = 87 else
"110111011111" when X = 30 AND Y = 87 else
"110111011111" when X = 31 AND Y = 87 else
"110111011111" when X = 32 AND Y = 87 else
"110111011111" when X = 33 AND Y = 87 else
"110111011111" when X = 34 AND Y = 87 else
"110111011111" when X = 35 AND Y = 87 else
"110111011111" when X = 36 AND Y = 87 else
"110111011111" when X = 37 AND Y = 87 else
"110111011111" when X = 38 AND Y = 87 else
"110111011111" when X = 39 AND Y = 87 else
"110111011111" when X = 40 AND Y = 87 else
"110111011111" when X = 41 AND Y = 87 else
"110111011111" when X = 42 AND Y = 87 else
"110111011111" when X = 43 AND Y = 87 else
"110111011111" when X = 44 AND Y = 87 else
"110111011111" when X = 45 AND Y = 87 else
"110111011111" when X = 46 AND Y = 87 else
"110111011111" when X = 47 AND Y = 87 else
"110111011111" when X = 48 AND Y = 87 else
"110111011111" when X = 49 AND Y = 87 else
"110111011111" when X = 50 AND Y = 87 else
"110111011111" when X = 51 AND Y = 87 else
"110111011111" when X = 52 AND Y = 87 else
"110111011111" when X = 53 AND Y = 87 else
"110111011111" when X = 54 AND Y = 87 else
"110111011111" when X = 55 AND Y = 87 else
"110111011111" when X = 56 AND Y = 87 else
"110111011111" when X = 57 AND Y = 87 else
"110111011111" when X = 58 AND Y = 87 else
"110111011111" when X = 59 AND Y = 87 else
"110111011111" when X = 60 AND Y = 87 else
"110111011111" when X = 61 AND Y = 87 else
"110111011111" when X = 62 AND Y = 87 else
"110111011111" when X = 63 AND Y = 87 else
"110111011111" when X = 64 AND Y = 87 else
"110111011111" when X = 65 AND Y = 87 else
"110111011111" when X = 66 AND Y = 87 else
"110111011111" when X = 67 AND Y = 87 else
"110111011111" when X = 68 AND Y = 87 else
"110111011111" when X = 69 AND Y = 87 else
"110111011111" when X = 70 AND Y = 87 else
"110111011111" when X = 71 AND Y = 87 else
"110111011111" when X = 72 AND Y = 87 else
"110111011111" when X = 73 AND Y = 87 else
"110111011111" when X = 74 AND Y = 87 else
"110111011111" when X = 75 AND Y = 87 else
"110111011111" when X = 76 AND Y = 87 else
"110111011111" when X = 77 AND Y = 87 else
"110111011111" when X = 78 AND Y = 87 else
"110111011111" when X = 79 AND Y = 87 else
"110111011111" when X = 80 AND Y = 87 else
"110111011111" when X = 81 AND Y = 87 else
"110111011111" when X = 82 AND Y = 87 else
"110111011111" when X = 83 AND Y = 87 else
"110111011111" when X = 84 AND Y = 87 else
"110111011111" when X = 85 AND Y = 87 else
"110111011111" when X = 86 AND Y = 87 else
"110111011111" when X = 87 AND Y = 87 else
"110111011111" when X = 88 AND Y = 87 else
"110111011111" when X = 89 AND Y = 87 else
"110111011111" when X = 90 AND Y = 87 else
"110111011111" when X = 91 AND Y = 87 else
"110111011111" when X = 92 AND Y = 87 else
"110111011111" when X = 93 AND Y = 87 else
"110111011111" when X = 94 AND Y = 87 else
"110111011111" when X = 95 AND Y = 87 else
"110111011111" when X = 96 AND Y = 87 else
"110111011111" when X = 97 AND Y = 87 else
"110111011111" when X = 98 AND Y = 87 else
"110111011111" when X = 99 AND Y = 87 else
"111111111111" when X = 100 AND Y = 87 else
"111111111111" when X = 101 AND Y = 87 else
"111111111111" when X = 102 AND Y = 87 else
"111111111111" when X = 103 AND Y = 87 else
"111111111111" when X = 104 AND Y = 87 else
"111111111111" when X = 105 AND Y = 87 else
"111111111111" when X = 106 AND Y = 87 else
"111111111111" when X = 107 AND Y = 87 else
"111111111111" when X = 108 AND Y = 87 else
"111111111111" when X = 109 AND Y = 87 else
"111111111111" when X = 110 AND Y = 87 else
"111111111111" when X = 111 AND Y = 87 else
"111111111111" when X = 112 AND Y = 87 else
"111111111111" when X = 113 AND Y = 87 else
"111111111111" when X = 114 AND Y = 87 else
"111111111111" when X = 115 AND Y = 87 else
"111111111111" when X = 116 AND Y = 87 else
"111111111111" when X = 117 AND Y = 87 else
"111111111111" when X = 118 AND Y = 87 else
"111111111111" when X = 119 AND Y = 87 else
"111111111111" when X = 120 AND Y = 87 else
"111111111111" when X = 121 AND Y = 87 else
"111111111111" when X = 122 AND Y = 87 else
"111111111111" when X = 123 AND Y = 87 else
"111111111111" when X = 124 AND Y = 87 else
"111111111111" when X = 125 AND Y = 87 else
"111111111111" when X = 126 AND Y = 87 else
"111111111111" when X = 127 AND Y = 87 else
"111111111111" when X = 128 AND Y = 87 else
"111111111111" when X = 129 AND Y = 87 else
"111111111111" when X = 130 AND Y = 87 else
"111111111111" when X = 131 AND Y = 87 else
"111111111111" when X = 132 AND Y = 87 else
"111111111111" when X = 133 AND Y = 87 else
"111111111111" when X = 134 AND Y = 87 else
"111111111111" when X = 135 AND Y = 87 else
"111111111111" when X = 136 AND Y = 87 else
"111111111111" when X = 137 AND Y = 87 else
"111111111111" when X = 138 AND Y = 87 else
"111111111111" when X = 139 AND Y = 87 else
"111111111111" when X = 140 AND Y = 87 else
"111111111111" when X = 141 AND Y = 87 else
"111111111111" when X = 142 AND Y = 87 else
"111111111111" when X = 143 AND Y = 87 else
"111111111111" when X = 144 AND Y = 87 else
"111111111111" when X = 145 AND Y = 87 else
"111111111111" when X = 146 AND Y = 87 else
"111111111111" when X = 147 AND Y = 87 else
"111111111111" when X = 148 AND Y = 87 else
"111111111111" when X = 149 AND Y = 87 else
"111111111111" when X = 150 AND Y = 87 else
"111111111111" when X = 151 AND Y = 87 else
"111111111111" when X = 152 AND Y = 87 else
"111111111111" when X = 153 AND Y = 87 else
"111111111111" when X = 154 AND Y = 87 else
"111111111111" when X = 155 AND Y = 87 else
"111111111111" when X = 156 AND Y = 87 else
"111111111111" when X = 157 AND Y = 87 else
"111111111111" when X = 158 AND Y = 87 else
"111111111111" when X = 159 AND Y = 87 else
"111111111111" when X = 160 AND Y = 87 else
"111111111111" when X = 161 AND Y = 87 else
"111111111111" when X = 162 AND Y = 87 else
"111111111111" when X = 163 AND Y = 87 else
"111111111111" when X = 164 AND Y = 87 else
"111111111111" when X = 165 AND Y = 87 else
"111111111111" when X = 166 AND Y = 87 else
"111111111111" when X = 167 AND Y = 87 else
"111111111111" when X = 168 AND Y = 87 else
"111111111111" when X = 169 AND Y = 87 else
"111111111111" when X = 170 AND Y = 87 else
"111111111111" when X = 171 AND Y = 87 else
"111111111111" when X = 172 AND Y = 87 else
"111111111111" when X = 173 AND Y = 87 else
"111111111111" when X = 174 AND Y = 87 else
"111111111111" when X = 175 AND Y = 87 else
"111111111111" when X = 176 AND Y = 87 else
"111111111111" when X = 177 AND Y = 87 else
"111111111111" when X = 178 AND Y = 87 else
"111111111111" when X = 179 AND Y = 87 else
"111111111111" when X = 180 AND Y = 87 else
"111111111111" when X = 181 AND Y = 87 else
"111111111111" when X = 182 AND Y = 87 else
"111111111111" when X = 183 AND Y = 87 else
"111111111111" when X = 184 AND Y = 87 else
"111111111111" when X = 185 AND Y = 87 else
"111111111111" when X = 186 AND Y = 87 else
"111111111111" when X = 187 AND Y = 87 else
"111111111111" when X = 188 AND Y = 87 else
"111111111111" when X = 189 AND Y = 87 else
"111111111111" when X = 190 AND Y = 87 else
"111111111111" when X = 191 AND Y = 87 else
"111111111111" when X = 192 AND Y = 87 else
"111111111111" when X = 193 AND Y = 87 else
"111111111111" when X = 194 AND Y = 87 else
"111111111111" when X = 195 AND Y = 87 else
"111111111111" when X = 196 AND Y = 87 else
"111111111111" when X = 197 AND Y = 87 else
"111111111111" when X = 198 AND Y = 87 else
"111111111111" when X = 199 AND Y = 87 else
"111111111111" when X = 200 AND Y = 87 else
"111111111111" when X = 201 AND Y = 87 else
"111111111111" when X = 202 AND Y = 87 else
"111111111111" when X = 203 AND Y = 87 else
"111111111111" when X = 204 AND Y = 87 else
"111111111111" when X = 205 AND Y = 87 else
"111111111111" when X = 206 AND Y = 87 else
"111111111111" when X = 207 AND Y = 87 else
"111111111111" when X = 208 AND Y = 87 else
"111111111111" when X = 209 AND Y = 87 else
"111111111111" when X = 210 AND Y = 87 else
"111111111111" when X = 211 AND Y = 87 else
"111111111111" when X = 212 AND Y = 87 else
"111111111111" when X = 213 AND Y = 87 else
"111111111111" when X = 214 AND Y = 87 else
"111111111111" when X = 215 AND Y = 87 else
"111111111111" when X = 216 AND Y = 87 else
"111111111111" when X = 217 AND Y = 87 else
"111111111111" when X = 218 AND Y = 87 else
"111111111111" when X = 219 AND Y = 87 else
"111111111111" when X = 220 AND Y = 87 else
"111111111111" when X = 221 AND Y = 87 else
"111111111111" when X = 222 AND Y = 87 else
"111111111111" when X = 223 AND Y = 87 else
"111111111111" when X = 224 AND Y = 87 else
"111111111111" when X = 225 AND Y = 87 else
"111111111111" when X = 226 AND Y = 87 else
"111111111111" when X = 227 AND Y = 87 else
"111111111111" when X = 228 AND Y = 87 else
"111111111111" when X = 229 AND Y = 87 else
"111111111111" when X = 230 AND Y = 87 else
"111111111111" when X = 231 AND Y = 87 else
"111111111111" when X = 232 AND Y = 87 else
"111111111111" when X = 233 AND Y = 87 else
"111111111111" when X = 234 AND Y = 87 else
"111111111111" when X = 235 AND Y = 87 else
"111111111111" when X = 236 AND Y = 87 else
"111111111111" when X = 237 AND Y = 87 else
"111111111111" when X = 238 AND Y = 87 else
"111111111111" when X = 239 AND Y = 87 else
"111111111111" when X = 240 AND Y = 87 else
"111111111111" when X = 241 AND Y = 87 else
"111111111111" when X = 242 AND Y = 87 else
"111111111111" when X = 243 AND Y = 87 else
"111111111111" when X = 244 AND Y = 87 else
"111111111111" when X = 245 AND Y = 87 else
"111111111111" when X = 246 AND Y = 87 else
"111111111111" when X = 247 AND Y = 87 else
"111111111111" when X = 248 AND Y = 87 else
"111111111111" when X = 249 AND Y = 87 else
"111111111111" when X = 250 AND Y = 87 else
"111111111111" when X = 251 AND Y = 87 else
"111111111111" when X = 252 AND Y = 87 else
"111111111111" when X = 253 AND Y = 87 else
"111111111111" when X = 254 AND Y = 87 else
"111111111111" when X = 255 AND Y = 87 else
"111111111111" when X = 256 AND Y = 87 else
"111111111111" when X = 257 AND Y = 87 else
"111111111111" when X = 258 AND Y = 87 else
"111111111111" when X = 259 AND Y = 87 else
"111111111111" when X = 260 AND Y = 87 else
"111111111111" when X = 261 AND Y = 87 else
"111111111111" when X = 262 AND Y = 87 else
"111111111111" when X = 263 AND Y = 87 else
"111111111111" when X = 264 AND Y = 87 else
"111111111111" when X = 265 AND Y = 87 else
"111111111111" when X = 266 AND Y = 87 else
"111111111111" when X = 267 AND Y = 87 else
"111111111111" when X = 268 AND Y = 87 else
"111111111111" when X = 269 AND Y = 87 else
"111111111111" when X = 270 AND Y = 87 else
"111111111111" when X = 271 AND Y = 87 else
"111111111111" when X = 272 AND Y = 87 else
"111111111111" when X = 273 AND Y = 87 else
"111111111111" when X = 274 AND Y = 87 else
"110111011111" when X = 275 AND Y = 87 else
"110111011111" when X = 276 AND Y = 87 else
"110111011111" when X = 277 AND Y = 87 else
"110111011111" when X = 278 AND Y = 87 else
"110111011111" when X = 279 AND Y = 87 else
"110111011111" when X = 280 AND Y = 87 else
"110111011111" when X = 281 AND Y = 87 else
"110111011111" when X = 282 AND Y = 87 else
"110111011111" when X = 283 AND Y = 87 else
"110111011111" when X = 284 AND Y = 87 else
"110111011111" when X = 285 AND Y = 87 else
"110111011111" when X = 286 AND Y = 87 else
"110111011111" when X = 287 AND Y = 87 else
"110111011111" when X = 288 AND Y = 87 else
"110111011111" when X = 289 AND Y = 87 else
"110111011111" when X = 290 AND Y = 87 else
"110111011111" when X = 291 AND Y = 87 else
"110111011111" when X = 292 AND Y = 87 else
"110111011111" when X = 293 AND Y = 87 else
"110111011111" when X = 294 AND Y = 87 else
"110111011111" when X = 295 AND Y = 87 else
"110111011111" when X = 296 AND Y = 87 else
"110111011111" when X = 297 AND Y = 87 else
"110111011111" when X = 298 AND Y = 87 else
"110111011111" when X = 299 AND Y = 87 else
"110111011111" when X = 300 AND Y = 87 else
"110111011111" when X = 301 AND Y = 87 else
"110111011111" when X = 302 AND Y = 87 else
"110111011111" when X = 303 AND Y = 87 else
"110111011111" when X = 304 AND Y = 87 else
"110111011111" when X = 305 AND Y = 87 else
"110111011111" when X = 306 AND Y = 87 else
"110111011111" when X = 307 AND Y = 87 else
"110111011111" when X = 308 AND Y = 87 else
"110111011111" when X = 309 AND Y = 87 else
"110111011111" when X = 310 AND Y = 87 else
"110111011111" when X = 311 AND Y = 87 else
"110111011111" when X = 312 AND Y = 87 else
"110111011111" when X = 313 AND Y = 87 else
"110111011111" when X = 314 AND Y = 87 else
"110111011111" when X = 315 AND Y = 87 else
"110111011111" when X = 316 AND Y = 87 else
"110111011111" when X = 317 AND Y = 87 else
"110111011111" when X = 318 AND Y = 87 else
"110111011111" when X = 319 AND Y = 87 else
"000000000000" when X = 320 AND Y = 87 else
"000000000000" when X = 321 AND Y = 87 else
"000000000000" when X = 322 AND Y = 87 else
"000000000000" when X = 323 AND Y = 87 else
"000000000000" when X = 324 AND Y = 87 else
"100010011101" when X = 0 AND Y = 88 else
"100010011101" when X = 1 AND Y = 88 else
"100010011101" when X = 2 AND Y = 88 else
"100010011101" when X = 3 AND Y = 88 else
"100010011101" when X = 4 AND Y = 88 else
"100010011101" when X = 5 AND Y = 88 else
"100010011101" when X = 6 AND Y = 88 else
"100010011101" when X = 7 AND Y = 88 else
"100010011101" when X = 8 AND Y = 88 else
"100010011101" when X = 9 AND Y = 88 else
"100010011101" when X = 10 AND Y = 88 else
"100010011101" when X = 11 AND Y = 88 else
"100010011101" when X = 12 AND Y = 88 else
"100010011101" when X = 13 AND Y = 88 else
"100010011101" when X = 14 AND Y = 88 else
"100010011101" when X = 15 AND Y = 88 else
"100010011101" when X = 16 AND Y = 88 else
"100010011101" when X = 17 AND Y = 88 else
"100010011101" when X = 18 AND Y = 88 else
"100010011101" when X = 19 AND Y = 88 else
"100010011101" when X = 20 AND Y = 88 else
"100010011101" when X = 21 AND Y = 88 else
"100010011101" when X = 22 AND Y = 88 else
"100010011101" when X = 23 AND Y = 88 else
"100010011101" when X = 24 AND Y = 88 else
"110111011111" when X = 25 AND Y = 88 else
"110111011111" when X = 26 AND Y = 88 else
"110111011111" when X = 27 AND Y = 88 else
"110111011111" when X = 28 AND Y = 88 else
"110111011111" when X = 29 AND Y = 88 else
"110111011111" when X = 30 AND Y = 88 else
"110111011111" when X = 31 AND Y = 88 else
"110111011111" when X = 32 AND Y = 88 else
"110111011111" when X = 33 AND Y = 88 else
"110111011111" when X = 34 AND Y = 88 else
"110111011111" when X = 35 AND Y = 88 else
"110111011111" when X = 36 AND Y = 88 else
"110111011111" when X = 37 AND Y = 88 else
"110111011111" when X = 38 AND Y = 88 else
"110111011111" when X = 39 AND Y = 88 else
"110111011111" when X = 40 AND Y = 88 else
"110111011111" when X = 41 AND Y = 88 else
"110111011111" when X = 42 AND Y = 88 else
"110111011111" when X = 43 AND Y = 88 else
"110111011111" when X = 44 AND Y = 88 else
"110111011111" when X = 45 AND Y = 88 else
"110111011111" when X = 46 AND Y = 88 else
"110111011111" when X = 47 AND Y = 88 else
"110111011111" when X = 48 AND Y = 88 else
"110111011111" when X = 49 AND Y = 88 else
"110111011111" when X = 50 AND Y = 88 else
"110111011111" when X = 51 AND Y = 88 else
"110111011111" when X = 52 AND Y = 88 else
"110111011111" when X = 53 AND Y = 88 else
"110111011111" when X = 54 AND Y = 88 else
"110111011111" when X = 55 AND Y = 88 else
"110111011111" when X = 56 AND Y = 88 else
"110111011111" when X = 57 AND Y = 88 else
"110111011111" when X = 58 AND Y = 88 else
"110111011111" when X = 59 AND Y = 88 else
"110111011111" when X = 60 AND Y = 88 else
"110111011111" when X = 61 AND Y = 88 else
"110111011111" when X = 62 AND Y = 88 else
"110111011111" when X = 63 AND Y = 88 else
"110111011111" when X = 64 AND Y = 88 else
"110111011111" when X = 65 AND Y = 88 else
"110111011111" when X = 66 AND Y = 88 else
"110111011111" when X = 67 AND Y = 88 else
"110111011111" when X = 68 AND Y = 88 else
"110111011111" when X = 69 AND Y = 88 else
"110111011111" when X = 70 AND Y = 88 else
"110111011111" when X = 71 AND Y = 88 else
"110111011111" when X = 72 AND Y = 88 else
"110111011111" when X = 73 AND Y = 88 else
"110111011111" when X = 74 AND Y = 88 else
"110111011111" when X = 75 AND Y = 88 else
"110111011111" when X = 76 AND Y = 88 else
"110111011111" when X = 77 AND Y = 88 else
"110111011111" when X = 78 AND Y = 88 else
"110111011111" when X = 79 AND Y = 88 else
"110111011111" when X = 80 AND Y = 88 else
"110111011111" when X = 81 AND Y = 88 else
"110111011111" when X = 82 AND Y = 88 else
"110111011111" when X = 83 AND Y = 88 else
"110111011111" when X = 84 AND Y = 88 else
"110111011111" when X = 85 AND Y = 88 else
"110111011111" when X = 86 AND Y = 88 else
"110111011111" when X = 87 AND Y = 88 else
"110111011111" when X = 88 AND Y = 88 else
"110111011111" when X = 89 AND Y = 88 else
"110111011111" when X = 90 AND Y = 88 else
"110111011111" when X = 91 AND Y = 88 else
"110111011111" when X = 92 AND Y = 88 else
"110111011111" when X = 93 AND Y = 88 else
"110111011111" when X = 94 AND Y = 88 else
"110111011111" when X = 95 AND Y = 88 else
"110111011111" when X = 96 AND Y = 88 else
"110111011111" when X = 97 AND Y = 88 else
"110111011111" when X = 98 AND Y = 88 else
"110111011111" when X = 99 AND Y = 88 else
"111111111111" when X = 100 AND Y = 88 else
"111111111111" when X = 101 AND Y = 88 else
"111111111111" when X = 102 AND Y = 88 else
"111111111111" when X = 103 AND Y = 88 else
"111111111111" when X = 104 AND Y = 88 else
"111111111111" when X = 105 AND Y = 88 else
"111111111111" when X = 106 AND Y = 88 else
"111111111111" when X = 107 AND Y = 88 else
"111111111111" when X = 108 AND Y = 88 else
"111111111111" when X = 109 AND Y = 88 else
"111111111111" when X = 110 AND Y = 88 else
"111111111111" when X = 111 AND Y = 88 else
"111111111111" when X = 112 AND Y = 88 else
"111111111111" when X = 113 AND Y = 88 else
"111111111111" when X = 114 AND Y = 88 else
"111111111111" when X = 115 AND Y = 88 else
"111111111111" when X = 116 AND Y = 88 else
"111111111111" when X = 117 AND Y = 88 else
"111111111111" when X = 118 AND Y = 88 else
"111111111111" when X = 119 AND Y = 88 else
"111111111111" when X = 120 AND Y = 88 else
"111111111111" when X = 121 AND Y = 88 else
"111111111111" when X = 122 AND Y = 88 else
"111111111111" when X = 123 AND Y = 88 else
"111111111111" when X = 124 AND Y = 88 else
"111111111111" when X = 125 AND Y = 88 else
"111111111111" when X = 126 AND Y = 88 else
"111111111111" when X = 127 AND Y = 88 else
"111111111111" when X = 128 AND Y = 88 else
"111111111111" when X = 129 AND Y = 88 else
"111111111111" when X = 130 AND Y = 88 else
"111111111111" when X = 131 AND Y = 88 else
"111111111111" when X = 132 AND Y = 88 else
"111111111111" when X = 133 AND Y = 88 else
"111111111111" when X = 134 AND Y = 88 else
"111111111111" when X = 135 AND Y = 88 else
"111111111111" when X = 136 AND Y = 88 else
"111111111111" when X = 137 AND Y = 88 else
"111111111111" when X = 138 AND Y = 88 else
"111111111111" when X = 139 AND Y = 88 else
"111111111111" when X = 140 AND Y = 88 else
"111111111111" when X = 141 AND Y = 88 else
"111111111111" when X = 142 AND Y = 88 else
"111111111111" when X = 143 AND Y = 88 else
"111111111111" when X = 144 AND Y = 88 else
"111111111111" when X = 145 AND Y = 88 else
"111111111111" when X = 146 AND Y = 88 else
"111111111111" when X = 147 AND Y = 88 else
"111111111111" when X = 148 AND Y = 88 else
"111111111111" when X = 149 AND Y = 88 else
"111111111111" when X = 150 AND Y = 88 else
"111111111111" when X = 151 AND Y = 88 else
"111111111111" when X = 152 AND Y = 88 else
"111111111111" when X = 153 AND Y = 88 else
"111111111111" when X = 154 AND Y = 88 else
"111111111111" when X = 155 AND Y = 88 else
"111111111111" when X = 156 AND Y = 88 else
"111111111111" when X = 157 AND Y = 88 else
"111111111111" when X = 158 AND Y = 88 else
"111111111111" when X = 159 AND Y = 88 else
"111111111111" when X = 160 AND Y = 88 else
"111111111111" when X = 161 AND Y = 88 else
"111111111111" when X = 162 AND Y = 88 else
"111111111111" when X = 163 AND Y = 88 else
"111111111111" when X = 164 AND Y = 88 else
"111111111111" when X = 165 AND Y = 88 else
"111111111111" when X = 166 AND Y = 88 else
"111111111111" when X = 167 AND Y = 88 else
"111111111111" when X = 168 AND Y = 88 else
"111111111111" when X = 169 AND Y = 88 else
"111111111111" when X = 170 AND Y = 88 else
"111111111111" when X = 171 AND Y = 88 else
"111111111111" when X = 172 AND Y = 88 else
"111111111111" when X = 173 AND Y = 88 else
"111111111111" when X = 174 AND Y = 88 else
"111111111111" when X = 175 AND Y = 88 else
"111111111111" when X = 176 AND Y = 88 else
"111111111111" when X = 177 AND Y = 88 else
"111111111111" when X = 178 AND Y = 88 else
"111111111111" when X = 179 AND Y = 88 else
"111111111111" when X = 180 AND Y = 88 else
"111111111111" when X = 181 AND Y = 88 else
"111111111111" when X = 182 AND Y = 88 else
"111111111111" when X = 183 AND Y = 88 else
"111111111111" when X = 184 AND Y = 88 else
"111111111111" when X = 185 AND Y = 88 else
"111111111111" when X = 186 AND Y = 88 else
"111111111111" when X = 187 AND Y = 88 else
"111111111111" when X = 188 AND Y = 88 else
"111111111111" when X = 189 AND Y = 88 else
"111111111111" when X = 190 AND Y = 88 else
"111111111111" when X = 191 AND Y = 88 else
"111111111111" when X = 192 AND Y = 88 else
"111111111111" when X = 193 AND Y = 88 else
"111111111111" when X = 194 AND Y = 88 else
"111111111111" when X = 195 AND Y = 88 else
"111111111111" when X = 196 AND Y = 88 else
"111111111111" when X = 197 AND Y = 88 else
"111111111111" when X = 198 AND Y = 88 else
"111111111111" when X = 199 AND Y = 88 else
"111111111111" when X = 200 AND Y = 88 else
"111111111111" when X = 201 AND Y = 88 else
"111111111111" when X = 202 AND Y = 88 else
"111111111111" when X = 203 AND Y = 88 else
"111111111111" when X = 204 AND Y = 88 else
"111111111111" when X = 205 AND Y = 88 else
"111111111111" when X = 206 AND Y = 88 else
"111111111111" when X = 207 AND Y = 88 else
"111111111111" when X = 208 AND Y = 88 else
"111111111111" when X = 209 AND Y = 88 else
"111111111111" when X = 210 AND Y = 88 else
"111111111111" when X = 211 AND Y = 88 else
"111111111111" when X = 212 AND Y = 88 else
"111111111111" when X = 213 AND Y = 88 else
"111111111111" when X = 214 AND Y = 88 else
"111111111111" when X = 215 AND Y = 88 else
"111111111111" when X = 216 AND Y = 88 else
"111111111111" when X = 217 AND Y = 88 else
"111111111111" when X = 218 AND Y = 88 else
"111111111111" when X = 219 AND Y = 88 else
"111111111111" when X = 220 AND Y = 88 else
"111111111111" when X = 221 AND Y = 88 else
"111111111111" when X = 222 AND Y = 88 else
"111111111111" when X = 223 AND Y = 88 else
"111111111111" when X = 224 AND Y = 88 else
"111111111111" when X = 225 AND Y = 88 else
"111111111111" when X = 226 AND Y = 88 else
"111111111111" when X = 227 AND Y = 88 else
"111111111111" when X = 228 AND Y = 88 else
"111111111111" when X = 229 AND Y = 88 else
"111111111111" when X = 230 AND Y = 88 else
"111111111111" when X = 231 AND Y = 88 else
"111111111111" when X = 232 AND Y = 88 else
"111111111111" when X = 233 AND Y = 88 else
"111111111111" when X = 234 AND Y = 88 else
"111111111111" when X = 235 AND Y = 88 else
"111111111111" when X = 236 AND Y = 88 else
"111111111111" when X = 237 AND Y = 88 else
"111111111111" when X = 238 AND Y = 88 else
"111111111111" when X = 239 AND Y = 88 else
"111111111111" when X = 240 AND Y = 88 else
"111111111111" when X = 241 AND Y = 88 else
"111111111111" when X = 242 AND Y = 88 else
"111111111111" when X = 243 AND Y = 88 else
"111111111111" when X = 244 AND Y = 88 else
"111111111111" when X = 245 AND Y = 88 else
"111111111111" when X = 246 AND Y = 88 else
"111111111111" when X = 247 AND Y = 88 else
"111111111111" when X = 248 AND Y = 88 else
"111111111111" when X = 249 AND Y = 88 else
"111111111111" when X = 250 AND Y = 88 else
"111111111111" when X = 251 AND Y = 88 else
"111111111111" when X = 252 AND Y = 88 else
"111111111111" when X = 253 AND Y = 88 else
"111111111111" when X = 254 AND Y = 88 else
"111111111111" when X = 255 AND Y = 88 else
"111111111111" when X = 256 AND Y = 88 else
"111111111111" when X = 257 AND Y = 88 else
"111111111111" when X = 258 AND Y = 88 else
"111111111111" when X = 259 AND Y = 88 else
"111111111111" when X = 260 AND Y = 88 else
"111111111111" when X = 261 AND Y = 88 else
"111111111111" when X = 262 AND Y = 88 else
"111111111111" when X = 263 AND Y = 88 else
"111111111111" when X = 264 AND Y = 88 else
"111111111111" when X = 265 AND Y = 88 else
"111111111111" when X = 266 AND Y = 88 else
"111111111111" when X = 267 AND Y = 88 else
"111111111111" when X = 268 AND Y = 88 else
"111111111111" when X = 269 AND Y = 88 else
"111111111111" when X = 270 AND Y = 88 else
"111111111111" when X = 271 AND Y = 88 else
"111111111111" when X = 272 AND Y = 88 else
"111111111111" when X = 273 AND Y = 88 else
"111111111111" when X = 274 AND Y = 88 else
"110111011111" when X = 275 AND Y = 88 else
"110111011111" when X = 276 AND Y = 88 else
"110111011111" when X = 277 AND Y = 88 else
"110111011111" when X = 278 AND Y = 88 else
"110111011111" when X = 279 AND Y = 88 else
"110111011111" when X = 280 AND Y = 88 else
"110111011111" when X = 281 AND Y = 88 else
"110111011111" when X = 282 AND Y = 88 else
"110111011111" when X = 283 AND Y = 88 else
"110111011111" when X = 284 AND Y = 88 else
"110111011111" when X = 285 AND Y = 88 else
"110111011111" when X = 286 AND Y = 88 else
"110111011111" when X = 287 AND Y = 88 else
"110111011111" when X = 288 AND Y = 88 else
"110111011111" when X = 289 AND Y = 88 else
"110111011111" when X = 290 AND Y = 88 else
"110111011111" when X = 291 AND Y = 88 else
"110111011111" when X = 292 AND Y = 88 else
"110111011111" when X = 293 AND Y = 88 else
"110111011111" when X = 294 AND Y = 88 else
"110111011111" when X = 295 AND Y = 88 else
"110111011111" when X = 296 AND Y = 88 else
"110111011111" when X = 297 AND Y = 88 else
"110111011111" when X = 298 AND Y = 88 else
"110111011111" when X = 299 AND Y = 88 else
"110111011111" when X = 300 AND Y = 88 else
"110111011111" when X = 301 AND Y = 88 else
"110111011111" when X = 302 AND Y = 88 else
"110111011111" when X = 303 AND Y = 88 else
"110111011111" when X = 304 AND Y = 88 else
"110111011111" when X = 305 AND Y = 88 else
"110111011111" when X = 306 AND Y = 88 else
"110111011111" when X = 307 AND Y = 88 else
"110111011111" when X = 308 AND Y = 88 else
"110111011111" when X = 309 AND Y = 88 else
"110111011111" when X = 310 AND Y = 88 else
"110111011111" when X = 311 AND Y = 88 else
"110111011111" when X = 312 AND Y = 88 else
"110111011111" when X = 313 AND Y = 88 else
"110111011111" when X = 314 AND Y = 88 else
"110111011111" when X = 315 AND Y = 88 else
"110111011111" when X = 316 AND Y = 88 else
"110111011111" when X = 317 AND Y = 88 else
"110111011111" when X = 318 AND Y = 88 else
"110111011111" when X = 319 AND Y = 88 else
"000000000000" when X = 320 AND Y = 88 else
"000000000000" when X = 321 AND Y = 88 else
"000000000000" when X = 322 AND Y = 88 else
"000000000000" when X = 323 AND Y = 88 else
"000000000000" when X = 324 AND Y = 88 else
"100010011101" when X = 0 AND Y = 89 else
"100010011101" when X = 1 AND Y = 89 else
"100010011101" when X = 2 AND Y = 89 else
"100010011101" when X = 3 AND Y = 89 else
"100010011101" when X = 4 AND Y = 89 else
"100010011101" when X = 5 AND Y = 89 else
"100010011101" when X = 6 AND Y = 89 else
"100010011101" when X = 7 AND Y = 89 else
"100010011101" when X = 8 AND Y = 89 else
"100010011101" when X = 9 AND Y = 89 else
"100010011101" when X = 10 AND Y = 89 else
"100010011101" when X = 11 AND Y = 89 else
"100010011101" when X = 12 AND Y = 89 else
"100010011101" when X = 13 AND Y = 89 else
"100010011101" when X = 14 AND Y = 89 else
"100010011101" when X = 15 AND Y = 89 else
"100010011101" when X = 16 AND Y = 89 else
"100010011101" when X = 17 AND Y = 89 else
"100010011101" when X = 18 AND Y = 89 else
"100010011101" when X = 19 AND Y = 89 else
"100010011101" when X = 20 AND Y = 89 else
"100010011101" when X = 21 AND Y = 89 else
"100010011101" when X = 22 AND Y = 89 else
"100010011101" when X = 23 AND Y = 89 else
"100010011101" when X = 24 AND Y = 89 else
"110111011111" when X = 25 AND Y = 89 else
"110111011111" when X = 26 AND Y = 89 else
"110111011111" when X = 27 AND Y = 89 else
"110111011111" when X = 28 AND Y = 89 else
"110111011111" when X = 29 AND Y = 89 else
"110111011111" when X = 30 AND Y = 89 else
"110111011111" when X = 31 AND Y = 89 else
"110111011111" when X = 32 AND Y = 89 else
"110111011111" when X = 33 AND Y = 89 else
"110111011111" when X = 34 AND Y = 89 else
"110111011111" when X = 35 AND Y = 89 else
"110111011111" when X = 36 AND Y = 89 else
"110111011111" when X = 37 AND Y = 89 else
"110111011111" when X = 38 AND Y = 89 else
"110111011111" when X = 39 AND Y = 89 else
"110111011111" when X = 40 AND Y = 89 else
"110111011111" when X = 41 AND Y = 89 else
"110111011111" when X = 42 AND Y = 89 else
"110111011111" when X = 43 AND Y = 89 else
"110111011111" when X = 44 AND Y = 89 else
"110111011111" when X = 45 AND Y = 89 else
"110111011111" when X = 46 AND Y = 89 else
"110111011111" when X = 47 AND Y = 89 else
"110111011111" when X = 48 AND Y = 89 else
"110111011111" when X = 49 AND Y = 89 else
"110111011111" when X = 50 AND Y = 89 else
"110111011111" when X = 51 AND Y = 89 else
"110111011111" when X = 52 AND Y = 89 else
"110111011111" when X = 53 AND Y = 89 else
"110111011111" when X = 54 AND Y = 89 else
"110111011111" when X = 55 AND Y = 89 else
"110111011111" when X = 56 AND Y = 89 else
"110111011111" when X = 57 AND Y = 89 else
"110111011111" when X = 58 AND Y = 89 else
"110111011111" when X = 59 AND Y = 89 else
"110111011111" when X = 60 AND Y = 89 else
"110111011111" when X = 61 AND Y = 89 else
"110111011111" when X = 62 AND Y = 89 else
"110111011111" when X = 63 AND Y = 89 else
"110111011111" when X = 64 AND Y = 89 else
"110111011111" when X = 65 AND Y = 89 else
"110111011111" when X = 66 AND Y = 89 else
"110111011111" when X = 67 AND Y = 89 else
"110111011111" when X = 68 AND Y = 89 else
"110111011111" when X = 69 AND Y = 89 else
"110111011111" when X = 70 AND Y = 89 else
"110111011111" when X = 71 AND Y = 89 else
"110111011111" when X = 72 AND Y = 89 else
"110111011111" when X = 73 AND Y = 89 else
"110111011111" when X = 74 AND Y = 89 else
"110111011111" when X = 75 AND Y = 89 else
"110111011111" when X = 76 AND Y = 89 else
"110111011111" when X = 77 AND Y = 89 else
"110111011111" when X = 78 AND Y = 89 else
"110111011111" when X = 79 AND Y = 89 else
"110111011111" when X = 80 AND Y = 89 else
"110111011111" when X = 81 AND Y = 89 else
"110111011111" when X = 82 AND Y = 89 else
"110111011111" when X = 83 AND Y = 89 else
"110111011111" when X = 84 AND Y = 89 else
"110111011111" when X = 85 AND Y = 89 else
"110111011111" when X = 86 AND Y = 89 else
"110111011111" when X = 87 AND Y = 89 else
"110111011111" when X = 88 AND Y = 89 else
"110111011111" when X = 89 AND Y = 89 else
"110111011111" when X = 90 AND Y = 89 else
"110111011111" when X = 91 AND Y = 89 else
"110111011111" when X = 92 AND Y = 89 else
"110111011111" when X = 93 AND Y = 89 else
"110111011111" when X = 94 AND Y = 89 else
"110111011111" when X = 95 AND Y = 89 else
"110111011111" when X = 96 AND Y = 89 else
"110111011111" when X = 97 AND Y = 89 else
"110111011111" when X = 98 AND Y = 89 else
"110111011111" when X = 99 AND Y = 89 else
"111111111111" when X = 100 AND Y = 89 else
"111111111111" when X = 101 AND Y = 89 else
"111111111111" when X = 102 AND Y = 89 else
"111111111111" when X = 103 AND Y = 89 else
"111111111111" when X = 104 AND Y = 89 else
"111111111111" when X = 105 AND Y = 89 else
"111111111111" when X = 106 AND Y = 89 else
"111111111111" when X = 107 AND Y = 89 else
"111111111111" when X = 108 AND Y = 89 else
"111111111111" when X = 109 AND Y = 89 else
"111111111111" when X = 110 AND Y = 89 else
"111111111111" when X = 111 AND Y = 89 else
"111111111111" when X = 112 AND Y = 89 else
"111111111111" when X = 113 AND Y = 89 else
"111111111111" when X = 114 AND Y = 89 else
"111111111111" when X = 115 AND Y = 89 else
"111111111111" when X = 116 AND Y = 89 else
"111111111111" when X = 117 AND Y = 89 else
"111111111111" when X = 118 AND Y = 89 else
"111111111111" when X = 119 AND Y = 89 else
"111111111111" when X = 120 AND Y = 89 else
"111111111111" when X = 121 AND Y = 89 else
"111111111111" when X = 122 AND Y = 89 else
"111111111111" when X = 123 AND Y = 89 else
"111111111111" when X = 124 AND Y = 89 else
"111111111111" when X = 125 AND Y = 89 else
"111111111111" when X = 126 AND Y = 89 else
"111111111111" when X = 127 AND Y = 89 else
"111111111111" when X = 128 AND Y = 89 else
"111111111111" when X = 129 AND Y = 89 else
"111111111111" when X = 130 AND Y = 89 else
"111111111111" when X = 131 AND Y = 89 else
"111111111111" when X = 132 AND Y = 89 else
"111111111111" when X = 133 AND Y = 89 else
"111111111111" when X = 134 AND Y = 89 else
"111111111111" when X = 135 AND Y = 89 else
"111111111111" when X = 136 AND Y = 89 else
"111111111111" when X = 137 AND Y = 89 else
"111111111111" when X = 138 AND Y = 89 else
"111111111111" when X = 139 AND Y = 89 else
"111111111111" when X = 140 AND Y = 89 else
"111111111111" when X = 141 AND Y = 89 else
"111111111111" when X = 142 AND Y = 89 else
"111111111111" when X = 143 AND Y = 89 else
"111111111111" when X = 144 AND Y = 89 else
"111111111111" when X = 145 AND Y = 89 else
"111111111111" when X = 146 AND Y = 89 else
"111111111111" when X = 147 AND Y = 89 else
"111111111111" when X = 148 AND Y = 89 else
"111111111111" when X = 149 AND Y = 89 else
"111111111111" when X = 150 AND Y = 89 else
"111111111111" when X = 151 AND Y = 89 else
"111111111111" when X = 152 AND Y = 89 else
"111111111111" when X = 153 AND Y = 89 else
"111111111111" when X = 154 AND Y = 89 else
"111111111111" when X = 155 AND Y = 89 else
"111111111111" when X = 156 AND Y = 89 else
"111111111111" when X = 157 AND Y = 89 else
"111111111111" when X = 158 AND Y = 89 else
"111111111111" when X = 159 AND Y = 89 else
"111111111111" when X = 160 AND Y = 89 else
"111111111111" when X = 161 AND Y = 89 else
"111111111111" when X = 162 AND Y = 89 else
"111111111111" when X = 163 AND Y = 89 else
"111111111111" when X = 164 AND Y = 89 else
"111111111111" when X = 165 AND Y = 89 else
"111111111111" when X = 166 AND Y = 89 else
"111111111111" when X = 167 AND Y = 89 else
"111111111111" when X = 168 AND Y = 89 else
"111111111111" when X = 169 AND Y = 89 else
"111111111111" when X = 170 AND Y = 89 else
"111111111111" when X = 171 AND Y = 89 else
"111111111111" when X = 172 AND Y = 89 else
"111111111111" when X = 173 AND Y = 89 else
"111111111111" when X = 174 AND Y = 89 else
"111111111111" when X = 175 AND Y = 89 else
"111111111111" when X = 176 AND Y = 89 else
"111111111111" when X = 177 AND Y = 89 else
"111111111111" when X = 178 AND Y = 89 else
"111111111111" when X = 179 AND Y = 89 else
"111111111111" when X = 180 AND Y = 89 else
"111111111111" when X = 181 AND Y = 89 else
"111111111111" when X = 182 AND Y = 89 else
"111111111111" when X = 183 AND Y = 89 else
"111111111111" when X = 184 AND Y = 89 else
"111111111111" when X = 185 AND Y = 89 else
"111111111111" when X = 186 AND Y = 89 else
"111111111111" when X = 187 AND Y = 89 else
"111111111111" when X = 188 AND Y = 89 else
"111111111111" when X = 189 AND Y = 89 else
"111111111111" when X = 190 AND Y = 89 else
"111111111111" when X = 191 AND Y = 89 else
"111111111111" when X = 192 AND Y = 89 else
"111111111111" when X = 193 AND Y = 89 else
"111111111111" when X = 194 AND Y = 89 else
"111111111111" when X = 195 AND Y = 89 else
"111111111111" when X = 196 AND Y = 89 else
"111111111111" when X = 197 AND Y = 89 else
"111111111111" when X = 198 AND Y = 89 else
"111111111111" when X = 199 AND Y = 89 else
"111111111111" when X = 200 AND Y = 89 else
"111111111111" when X = 201 AND Y = 89 else
"111111111111" when X = 202 AND Y = 89 else
"111111111111" when X = 203 AND Y = 89 else
"111111111111" when X = 204 AND Y = 89 else
"111111111111" when X = 205 AND Y = 89 else
"111111111111" when X = 206 AND Y = 89 else
"111111111111" when X = 207 AND Y = 89 else
"111111111111" when X = 208 AND Y = 89 else
"111111111111" when X = 209 AND Y = 89 else
"111111111111" when X = 210 AND Y = 89 else
"111111111111" when X = 211 AND Y = 89 else
"111111111111" when X = 212 AND Y = 89 else
"111111111111" when X = 213 AND Y = 89 else
"111111111111" when X = 214 AND Y = 89 else
"111111111111" when X = 215 AND Y = 89 else
"111111111111" when X = 216 AND Y = 89 else
"111111111111" when X = 217 AND Y = 89 else
"111111111111" when X = 218 AND Y = 89 else
"111111111111" when X = 219 AND Y = 89 else
"111111111111" when X = 220 AND Y = 89 else
"111111111111" when X = 221 AND Y = 89 else
"111111111111" when X = 222 AND Y = 89 else
"111111111111" when X = 223 AND Y = 89 else
"111111111111" when X = 224 AND Y = 89 else
"111111111111" when X = 225 AND Y = 89 else
"111111111111" when X = 226 AND Y = 89 else
"111111111111" when X = 227 AND Y = 89 else
"111111111111" when X = 228 AND Y = 89 else
"111111111111" when X = 229 AND Y = 89 else
"111111111111" when X = 230 AND Y = 89 else
"111111111111" when X = 231 AND Y = 89 else
"111111111111" when X = 232 AND Y = 89 else
"111111111111" when X = 233 AND Y = 89 else
"111111111111" when X = 234 AND Y = 89 else
"111111111111" when X = 235 AND Y = 89 else
"111111111111" when X = 236 AND Y = 89 else
"111111111111" when X = 237 AND Y = 89 else
"111111111111" when X = 238 AND Y = 89 else
"111111111111" when X = 239 AND Y = 89 else
"111111111111" when X = 240 AND Y = 89 else
"111111111111" when X = 241 AND Y = 89 else
"111111111111" when X = 242 AND Y = 89 else
"111111111111" when X = 243 AND Y = 89 else
"111111111111" when X = 244 AND Y = 89 else
"111111111111" when X = 245 AND Y = 89 else
"111111111111" when X = 246 AND Y = 89 else
"111111111111" when X = 247 AND Y = 89 else
"111111111111" when X = 248 AND Y = 89 else
"111111111111" when X = 249 AND Y = 89 else
"111111111111" when X = 250 AND Y = 89 else
"111111111111" when X = 251 AND Y = 89 else
"111111111111" when X = 252 AND Y = 89 else
"111111111111" when X = 253 AND Y = 89 else
"111111111111" when X = 254 AND Y = 89 else
"111111111111" when X = 255 AND Y = 89 else
"111111111111" when X = 256 AND Y = 89 else
"111111111111" when X = 257 AND Y = 89 else
"111111111111" when X = 258 AND Y = 89 else
"111111111111" when X = 259 AND Y = 89 else
"111111111111" when X = 260 AND Y = 89 else
"111111111111" when X = 261 AND Y = 89 else
"111111111111" when X = 262 AND Y = 89 else
"111111111111" when X = 263 AND Y = 89 else
"111111111111" when X = 264 AND Y = 89 else
"111111111111" when X = 265 AND Y = 89 else
"111111111111" when X = 266 AND Y = 89 else
"111111111111" when X = 267 AND Y = 89 else
"111111111111" when X = 268 AND Y = 89 else
"111111111111" when X = 269 AND Y = 89 else
"111111111111" when X = 270 AND Y = 89 else
"111111111111" when X = 271 AND Y = 89 else
"111111111111" when X = 272 AND Y = 89 else
"111111111111" when X = 273 AND Y = 89 else
"111111111111" when X = 274 AND Y = 89 else
"110111011111" when X = 275 AND Y = 89 else
"110111011111" when X = 276 AND Y = 89 else
"110111011111" when X = 277 AND Y = 89 else
"110111011111" when X = 278 AND Y = 89 else
"110111011111" when X = 279 AND Y = 89 else
"110111011111" when X = 280 AND Y = 89 else
"110111011111" when X = 281 AND Y = 89 else
"110111011111" when X = 282 AND Y = 89 else
"110111011111" when X = 283 AND Y = 89 else
"110111011111" when X = 284 AND Y = 89 else
"110111011111" when X = 285 AND Y = 89 else
"110111011111" when X = 286 AND Y = 89 else
"110111011111" when X = 287 AND Y = 89 else
"110111011111" when X = 288 AND Y = 89 else
"110111011111" when X = 289 AND Y = 89 else
"110111011111" when X = 290 AND Y = 89 else
"110111011111" when X = 291 AND Y = 89 else
"110111011111" when X = 292 AND Y = 89 else
"110111011111" when X = 293 AND Y = 89 else
"110111011111" when X = 294 AND Y = 89 else
"110111011111" when X = 295 AND Y = 89 else
"110111011111" when X = 296 AND Y = 89 else
"110111011111" when X = 297 AND Y = 89 else
"110111011111" when X = 298 AND Y = 89 else
"110111011111" when X = 299 AND Y = 89 else
"110111011111" when X = 300 AND Y = 89 else
"110111011111" when X = 301 AND Y = 89 else
"110111011111" when X = 302 AND Y = 89 else
"110111011111" when X = 303 AND Y = 89 else
"110111011111" when X = 304 AND Y = 89 else
"110111011111" when X = 305 AND Y = 89 else
"110111011111" when X = 306 AND Y = 89 else
"110111011111" when X = 307 AND Y = 89 else
"110111011111" when X = 308 AND Y = 89 else
"110111011111" when X = 309 AND Y = 89 else
"110111011111" when X = 310 AND Y = 89 else
"110111011111" when X = 311 AND Y = 89 else
"110111011111" when X = 312 AND Y = 89 else
"110111011111" when X = 313 AND Y = 89 else
"110111011111" when X = 314 AND Y = 89 else
"110111011111" when X = 315 AND Y = 89 else
"110111011111" when X = 316 AND Y = 89 else
"110111011111" when X = 317 AND Y = 89 else
"110111011111" when X = 318 AND Y = 89 else
"110111011111" when X = 319 AND Y = 89 else
"000000000000" when X = 320 AND Y = 89 else
"000000000000" when X = 321 AND Y = 89 else
"000000000000" when X = 322 AND Y = 89 else
"000000000000" when X = 323 AND Y = 89 else
"000000000000" when X = 324 AND Y = 89 else
"100010011101" when X = 0 AND Y = 90 else
"100010011101" when X = 1 AND Y = 90 else
"100010011101" when X = 2 AND Y = 90 else
"100010011101" when X = 3 AND Y = 90 else
"100010011101" when X = 4 AND Y = 90 else
"100010011101" when X = 5 AND Y = 90 else
"100010011101" when X = 6 AND Y = 90 else
"100010011101" when X = 7 AND Y = 90 else
"100010011101" when X = 8 AND Y = 90 else
"100010011101" when X = 9 AND Y = 90 else
"100010011101" when X = 10 AND Y = 90 else
"100010011101" when X = 11 AND Y = 90 else
"100010011101" when X = 12 AND Y = 90 else
"100010011101" when X = 13 AND Y = 90 else
"100010011101" when X = 14 AND Y = 90 else
"100010011101" when X = 15 AND Y = 90 else
"100010011101" when X = 16 AND Y = 90 else
"100010011101" when X = 17 AND Y = 90 else
"100010011101" when X = 18 AND Y = 90 else
"100010011101" when X = 19 AND Y = 90 else
"110111011111" when X = 20 AND Y = 90 else
"110111011111" when X = 21 AND Y = 90 else
"110111011111" when X = 22 AND Y = 90 else
"110111011111" when X = 23 AND Y = 90 else
"110111011111" when X = 24 AND Y = 90 else
"110111011111" when X = 25 AND Y = 90 else
"110111011111" when X = 26 AND Y = 90 else
"110111011111" when X = 27 AND Y = 90 else
"110111011111" when X = 28 AND Y = 90 else
"110111011111" when X = 29 AND Y = 90 else
"110111011111" when X = 30 AND Y = 90 else
"110111011111" when X = 31 AND Y = 90 else
"110111011111" when X = 32 AND Y = 90 else
"110111011111" when X = 33 AND Y = 90 else
"110111011111" when X = 34 AND Y = 90 else
"110111011111" when X = 35 AND Y = 90 else
"110111011111" when X = 36 AND Y = 90 else
"110111011111" when X = 37 AND Y = 90 else
"110111011111" when X = 38 AND Y = 90 else
"110111011111" when X = 39 AND Y = 90 else
"110111011111" when X = 40 AND Y = 90 else
"110111011111" when X = 41 AND Y = 90 else
"110111011111" when X = 42 AND Y = 90 else
"110111011111" when X = 43 AND Y = 90 else
"110111011111" when X = 44 AND Y = 90 else
"110111011111" when X = 45 AND Y = 90 else
"110111011111" when X = 46 AND Y = 90 else
"110111011111" when X = 47 AND Y = 90 else
"110111011111" when X = 48 AND Y = 90 else
"110111011111" when X = 49 AND Y = 90 else
"110111011111" when X = 50 AND Y = 90 else
"110111011111" when X = 51 AND Y = 90 else
"110111011111" when X = 52 AND Y = 90 else
"110111011111" when X = 53 AND Y = 90 else
"110111011111" when X = 54 AND Y = 90 else
"110111011111" when X = 55 AND Y = 90 else
"110111011111" when X = 56 AND Y = 90 else
"110111011111" when X = 57 AND Y = 90 else
"110111011111" when X = 58 AND Y = 90 else
"110111011111" when X = 59 AND Y = 90 else
"110111011111" when X = 60 AND Y = 90 else
"110111011111" when X = 61 AND Y = 90 else
"110111011111" when X = 62 AND Y = 90 else
"110111011111" when X = 63 AND Y = 90 else
"110111011111" when X = 64 AND Y = 90 else
"110111011111" when X = 65 AND Y = 90 else
"110111011111" when X = 66 AND Y = 90 else
"110111011111" when X = 67 AND Y = 90 else
"110111011111" when X = 68 AND Y = 90 else
"110111011111" when X = 69 AND Y = 90 else
"111111111111" when X = 70 AND Y = 90 else
"111111111111" when X = 71 AND Y = 90 else
"111111111111" when X = 72 AND Y = 90 else
"111111111111" when X = 73 AND Y = 90 else
"111111111111" when X = 74 AND Y = 90 else
"111111111111" when X = 75 AND Y = 90 else
"111111111111" when X = 76 AND Y = 90 else
"111111111111" when X = 77 AND Y = 90 else
"111111111111" when X = 78 AND Y = 90 else
"111111111111" when X = 79 AND Y = 90 else
"111111111111" when X = 80 AND Y = 90 else
"111111111111" when X = 81 AND Y = 90 else
"111111111111" when X = 82 AND Y = 90 else
"111111111111" when X = 83 AND Y = 90 else
"111111111111" when X = 84 AND Y = 90 else
"111111111111" when X = 85 AND Y = 90 else
"111111111111" when X = 86 AND Y = 90 else
"111111111111" when X = 87 AND Y = 90 else
"111111111111" when X = 88 AND Y = 90 else
"111111111111" when X = 89 AND Y = 90 else
"111111111111" when X = 90 AND Y = 90 else
"111111111111" when X = 91 AND Y = 90 else
"111111111111" when X = 92 AND Y = 90 else
"111111111111" when X = 93 AND Y = 90 else
"111111111111" when X = 94 AND Y = 90 else
"111111111111" when X = 95 AND Y = 90 else
"111111111111" when X = 96 AND Y = 90 else
"111111111111" when X = 97 AND Y = 90 else
"111111111111" when X = 98 AND Y = 90 else
"111111111111" when X = 99 AND Y = 90 else
"111111111111" when X = 100 AND Y = 90 else
"111111111111" when X = 101 AND Y = 90 else
"111111111111" when X = 102 AND Y = 90 else
"111111111111" when X = 103 AND Y = 90 else
"111111111111" when X = 104 AND Y = 90 else
"111111111111" when X = 105 AND Y = 90 else
"111111111111" when X = 106 AND Y = 90 else
"111111111111" when X = 107 AND Y = 90 else
"111111111111" when X = 108 AND Y = 90 else
"111111111111" when X = 109 AND Y = 90 else
"111111111111" when X = 110 AND Y = 90 else
"111111111111" when X = 111 AND Y = 90 else
"111111111111" when X = 112 AND Y = 90 else
"111111111111" when X = 113 AND Y = 90 else
"111111111111" when X = 114 AND Y = 90 else
"111111111111" when X = 115 AND Y = 90 else
"111111111111" when X = 116 AND Y = 90 else
"111111111111" when X = 117 AND Y = 90 else
"111111111111" when X = 118 AND Y = 90 else
"111111111111" when X = 119 AND Y = 90 else
"111111111111" when X = 120 AND Y = 90 else
"111111111111" when X = 121 AND Y = 90 else
"111111111111" when X = 122 AND Y = 90 else
"111111111111" when X = 123 AND Y = 90 else
"111111111111" when X = 124 AND Y = 90 else
"111111111111" when X = 125 AND Y = 90 else
"111111111111" when X = 126 AND Y = 90 else
"111111111111" when X = 127 AND Y = 90 else
"111111111111" when X = 128 AND Y = 90 else
"111111111111" when X = 129 AND Y = 90 else
"111111111111" when X = 130 AND Y = 90 else
"111111111111" when X = 131 AND Y = 90 else
"111111111111" when X = 132 AND Y = 90 else
"111111111111" when X = 133 AND Y = 90 else
"111111111111" when X = 134 AND Y = 90 else
"111111111111" when X = 135 AND Y = 90 else
"111111111111" when X = 136 AND Y = 90 else
"111111111111" when X = 137 AND Y = 90 else
"111111111111" when X = 138 AND Y = 90 else
"111111111111" when X = 139 AND Y = 90 else
"111111111111" when X = 140 AND Y = 90 else
"111111111111" when X = 141 AND Y = 90 else
"111111111111" when X = 142 AND Y = 90 else
"111111111111" when X = 143 AND Y = 90 else
"111111111111" when X = 144 AND Y = 90 else
"111111111111" when X = 145 AND Y = 90 else
"111111111111" when X = 146 AND Y = 90 else
"111111111111" when X = 147 AND Y = 90 else
"111111111111" when X = 148 AND Y = 90 else
"111111111111" when X = 149 AND Y = 90 else
"111111111111" when X = 150 AND Y = 90 else
"111111111111" when X = 151 AND Y = 90 else
"111111111111" when X = 152 AND Y = 90 else
"111111111111" when X = 153 AND Y = 90 else
"111111111111" when X = 154 AND Y = 90 else
"111111111111" when X = 155 AND Y = 90 else
"111111111111" when X = 156 AND Y = 90 else
"111111111111" when X = 157 AND Y = 90 else
"111111111111" when X = 158 AND Y = 90 else
"111111111111" when X = 159 AND Y = 90 else
"111111111111" when X = 160 AND Y = 90 else
"111111111111" when X = 161 AND Y = 90 else
"111111111111" when X = 162 AND Y = 90 else
"111111111111" when X = 163 AND Y = 90 else
"111111111111" when X = 164 AND Y = 90 else
"111111111111" when X = 165 AND Y = 90 else
"111111111111" when X = 166 AND Y = 90 else
"111111111111" when X = 167 AND Y = 90 else
"111111111111" when X = 168 AND Y = 90 else
"111111111111" when X = 169 AND Y = 90 else
"111111111111" when X = 170 AND Y = 90 else
"111111111111" when X = 171 AND Y = 90 else
"111111111111" when X = 172 AND Y = 90 else
"111111111111" when X = 173 AND Y = 90 else
"111111111111" when X = 174 AND Y = 90 else
"111111111111" when X = 175 AND Y = 90 else
"111111111111" when X = 176 AND Y = 90 else
"111111111111" when X = 177 AND Y = 90 else
"111111111111" when X = 178 AND Y = 90 else
"111111111111" when X = 179 AND Y = 90 else
"111111111111" when X = 180 AND Y = 90 else
"111111111111" when X = 181 AND Y = 90 else
"111111111111" when X = 182 AND Y = 90 else
"111111111111" when X = 183 AND Y = 90 else
"111111111111" when X = 184 AND Y = 90 else
"111111111111" when X = 185 AND Y = 90 else
"111111111111" when X = 186 AND Y = 90 else
"111111111111" when X = 187 AND Y = 90 else
"111111111111" when X = 188 AND Y = 90 else
"111111111111" when X = 189 AND Y = 90 else
"111111111111" when X = 190 AND Y = 90 else
"111111111111" when X = 191 AND Y = 90 else
"111111111111" when X = 192 AND Y = 90 else
"111111111111" when X = 193 AND Y = 90 else
"111111111111" when X = 194 AND Y = 90 else
"111111111111" when X = 195 AND Y = 90 else
"111111111111" when X = 196 AND Y = 90 else
"111111111111" when X = 197 AND Y = 90 else
"111111111111" when X = 198 AND Y = 90 else
"111111111111" when X = 199 AND Y = 90 else
"111111111111" when X = 200 AND Y = 90 else
"111111111111" when X = 201 AND Y = 90 else
"111111111111" when X = 202 AND Y = 90 else
"111111111111" when X = 203 AND Y = 90 else
"111111111111" when X = 204 AND Y = 90 else
"111111111111" when X = 205 AND Y = 90 else
"111111111111" when X = 206 AND Y = 90 else
"111111111111" when X = 207 AND Y = 90 else
"111111111111" when X = 208 AND Y = 90 else
"111111111111" when X = 209 AND Y = 90 else
"111111111111" when X = 210 AND Y = 90 else
"111111111111" when X = 211 AND Y = 90 else
"111111111111" when X = 212 AND Y = 90 else
"111111111111" when X = 213 AND Y = 90 else
"111111111111" when X = 214 AND Y = 90 else
"111111111111" when X = 215 AND Y = 90 else
"111111111111" when X = 216 AND Y = 90 else
"111111111111" when X = 217 AND Y = 90 else
"111111111111" when X = 218 AND Y = 90 else
"111111111111" when X = 219 AND Y = 90 else
"110111011111" when X = 220 AND Y = 90 else
"110111011111" when X = 221 AND Y = 90 else
"110111011111" when X = 222 AND Y = 90 else
"110111011111" when X = 223 AND Y = 90 else
"110111011111" when X = 224 AND Y = 90 else
"110111011111" when X = 225 AND Y = 90 else
"110111011111" when X = 226 AND Y = 90 else
"110111011111" when X = 227 AND Y = 90 else
"110111011111" when X = 228 AND Y = 90 else
"110111011111" when X = 229 AND Y = 90 else
"111111111111" when X = 230 AND Y = 90 else
"111111111111" when X = 231 AND Y = 90 else
"111111111111" when X = 232 AND Y = 90 else
"111111111111" when X = 233 AND Y = 90 else
"111111111111" when X = 234 AND Y = 90 else
"111111111111" when X = 235 AND Y = 90 else
"111111111111" when X = 236 AND Y = 90 else
"111111111111" when X = 237 AND Y = 90 else
"111111111111" when X = 238 AND Y = 90 else
"111111111111" when X = 239 AND Y = 90 else
"111111111111" when X = 240 AND Y = 90 else
"111111111111" when X = 241 AND Y = 90 else
"111111111111" when X = 242 AND Y = 90 else
"111111111111" when X = 243 AND Y = 90 else
"111111111111" when X = 244 AND Y = 90 else
"111111111111" when X = 245 AND Y = 90 else
"111111111111" when X = 246 AND Y = 90 else
"111111111111" when X = 247 AND Y = 90 else
"111111111111" when X = 248 AND Y = 90 else
"111111111111" when X = 249 AND Y = 90 else
"111111111111" when X = 250 AND Y = 90 else
"111111111111" when X = 251 AND Y = 90 else
"111111111111" when X = 252 AND Y = 90 else
"111111111111" when X = 253 AND Y = 90 else
"111111111111" when X = 254 AND Y = 90 else
"111111111111" when X = 255 AND Y = 90 else
"111111111111" when X = 256 AND Y = 90 else
"111111111111" when X = 257 AND Y = 90 else
"111111111111" when X = 258 AND Y = 90 else
"111111111111" when X = 259 AND Y = 90 else
"111111111111" when X = 260 AND Y = 90 else
"111111111111" when X = 261 AND Y = 90 else
"111111111111" when X = 262 AND Y = 90 else
"111111111111" when X = 263 AND Y = 90 else
"111111111111" when X = 264 AND Y = 90 else
"111111111111" when X = 265 AND Y = 90 else
"111111111111" when X = 266 AND Y = 90 else
"111111111111" when X = 267 AND Y = 90 else
"111111111111" when X = 268 AND Y = 90 else
"111111111111" when X = 269 AND Y = 90 else
"111111111111" when X = 270 AND Y = 90 else
"111111111111" when X = 271 AND Y = 90 else
"111111111111" when X = 272 AND Y = 90 else
"111111111111" when X = 273 AND Y = 90 else
"111111111111" when X = 274 AND Y = 90 else
"110111011111" when X = 275 AND Y = 90 else
"110111011111" when X = 276 AND Y = 90 else
"110111011111" when X = 277 AND Y = 90 else
"110111011111" when X = 278 AND Y = 90 else
"110111011111" when X = 279 AND Y = 90 else
"110111011111" when X = 280 AND Y = 90 else
"110111011111" when X = 281 AND Y = 90 else
"110111011111" when X = 282 AND Y = 90 else
"110111011111" when X = 283 AND Y = 90 else
"110111011111" when X = 284 AND Y = 90 else
"110111011111" when X = 285 AND Y = 90 else
"110111011111" when X = 286 AND Y = 90 else
"110111011111" when X = 287 AND Y = 90 else
"110111011111" when X = 288 AND Y = 90 else
"110111011111" when X = 289 AND Y = 90 else
"110111011111" when X = 290 AND Y = 90 else
"110111011111" when X = 291 AND Y = 90 else
"110111011111" when X = 292 AND Y = 90 else
"110111011111" when X = 293 AND Y = 90 else
"110111011111" when X = 294 AND Y = 90 else
"110111011111" when X = 295 AND Y = 90 else
"110111011111" when X = 296 AND Y = 90 else
"110111011111" when X = 297 AND Y = 90 else
"110111011111" when X = 298 AND Y = 90 else
"110111011111" when X = 299 AND Y = 90 else
"110111011111" when X = 300 AND Y = 90 else
"110111011111" when X = 301 AND Y = 90 else
"110111011111" when X = 302 AND Y = 90 else
"110111011111" when X = 303 AND Y = 90 else
"110111011111" when X = 304 AND Y = 90 else
"110111011111" when X = 305 AND Y = 90 else
"110111011111" when X = 306 AND Y = 90 else
"110111011111" when X = 307 AND Y = 90 else
"110111011111" when X = 308 AND Y = 90 else
"110111011111" when X = 309 AND Y = 90 else
"110111011111" when X = 310 AND Y = 90 else
"110111011111" when X = 311 AND Y = 90 else
"110111011111" when X = 312 AND Y = 90 else
"110111011111" when X = 313 AND Y = 90 else
"110111011111" when X = 314 AND Y = 90 else
"110111011111" when X = 315 AND Y = 90 else
"110111011111" when X = 316 AND Y = 90 else
"110111011111" when X = 317 AND Y = 90 else
"110111011111" when X = 318 AND Y = 90 else
"110111011111" when X = 319 AND Y = 90 else
"000000000000" when X = 320 AND Y = 90 else
"000000000000" when X = 321 AND Y = 90 else
"000000000000" when X = 322 AND Y = 90 else
"000000000000" when X = 323 AND Y = 90 else
"000000000000" when X = 324 AND Y = 90 else
"100010011101" when X = 0 AND Y = 91 else
"100010011101" when X = 1 AND Y = 91 else
"100010011101" when X = 2 AND Y = 91 else
"100010011101" when X = 3 AND Y = 91 else
"100010011101" when X = 4 AND Y = 91 else
"100010011101" when X = 5 AND Y = 91 else
"100010011101" when X = 6 AND Y = 91 else
"100010011101" when X = 7 AND Y = 91 else
"100010011101" when X = 8 AND Y = 91 else
"100010011101" when X = 9 AND Y = 91 else
"100010011101" when X = 10 AND Y = 91 else
"100010011101" when X = 11 AND Y = 91 else
"100010011101" when X = 12 AND Y = 91 else
"100010011101" when X = 13 AND Y = 91 else
"100010011101" when X = 14 AND Y = 91 else
"100010011101" when X = 15 AND Y = 91 else
"100010011101" when X = 16 AND Y = 91 else
"100010011101" when X = 17 AND Y = 91 else
"100010011101" when X = 18 AND Y = 91 else
"100010011101" when X = 19 AND Y = 91 else
"110111011111" when X = 20 AND Y = 91 else
"110111011111" when X = 21 AND Y = 91 else
"110111011111" when X = 22 AND Y = 91 else
"110111011111" when X = 23 AND Y = 91 else
"110111011111" when X = 24 AND Y = 91 else
"110111011111" when X = 25 AND Y = 91 else
"110111011111" when X = 26 AND Y = 91 else
"110111011111" when X = 27 AND Y = 91 else
"110111011111" when X = 28 AND Y = 91 else
"110111011111" when X = 29 AND Y = 91 else
"110111011111" when X = 30 AND Y = 91 else
"110111011111" when X = 31 AND Y = 91 else
"110111011111" when X = 32 AND Y = 91 else
"110111011111" when X = 33 AND Y = 91 else
"110111011111" when X = 34 AND Y = 91 else
"110111011111" when X = 35 AND Y = 91 else
"110111011111" when X = 36 AND Y = 91 else
"110111011111" when X = 37 AND Y = 91 else
"110111011111" when X = 38 AND Y = 91 else
"110111011111" when X = 39 AND Y = 91 else
"110111011111" when X = 40 AND Y = 91 else
"110111011111" when X = 41 AND Y = 91 else
"110111011111" when X = 42 AND Y = 91 else
"110111011111" when X = 43 AND Y = 91 else
"110111011111" when X = 44 AND Y = 91 else
"110111011111" when X = 45 AND Y = 91 else
"110111011111" when X = 46 AND Y = 91 else
"110111011111" when X = 47 AND Y = 91 else
"110111011111" when X = 48 AND Y = 91 else
"110111011111" when X = 49 AND Y = 91 else
"110111011111" when X = 50 AND Y = 91 else
"110111011111" when X = 51 AND Y = 91 else
"110111011111" when X = 52 AND Y = 91 else
"110111011111" when X = 53 AND Y = 91 else
"110111011111" when X = 54 AND Y = 91 else
"110111011111" when X = 55 AND Y = 91 else
"110111011111" when X = 56 AND Y = 91 else
"110111011111" when X = 57 AND Y = 91 else
"110111011111" when X = 58 AND Y = 91 else
"110111011111" when X = 59 AND Y = 91 else
"110111011111" when X = 60 AND Y = 91 else
"110111011111" when X = 61 AND Y = 91 else
"110111011111" when X = 62 AND Y = 91 else
"110111011111" when X = 63 AND Y = 91 else
"110111011111" when X = 64 AND Y = 91 else
"110111011111" when X = 65 AND Y = 91 else
"110111011111" when X = 66 AND Y = 91 else
"110111011111" when X = 67 AND Y = 91 else
"110111011111" when X = 68 AND Y = 91 else
"110111011111" when X = 69 AND Y = 91 else
"111111111111" when X = 70 AND Y = 91 else
"111111111111" when X = 71 AND Y = 91 else
"111111111111" when X = 72 AND Y = 91 else
"111111111111" when X = 73 AND Y = 91 else
"111111111111" when X = 74 AND Y = 91 else
"111111111111" when X = 75 AND Y = 91 else
"111111111111" when X = 76 AND Y = 91 else
"111111111111" when X = 77 AND Y = 91 else
"111111111111" when X = 78 AND Y = 91 else
"111111111111" when X = 79 AND Y = 91 else
"111111111111" when X = 80 AND Y = 91 else
"111111111111" when X = 81 AND Y = 91 else
"111111111111" when X = 82 AND Y = 91 else
"111111111111" when X = 83 AND Y = 91 else
"111111111111" when X = 84 AND Y = 91 else
"111111111111" when X = 85 AND Y = 91 else
"111111111111" when X = 86 AND Y = 91 else
"111111111111" when X = 87 AND Y = 91 else
"111111111111" when X = 88 AND Y = 91 else
"111111111111" when X = 89 AND Y = 91 else
"111111111111" when X = 90 AND Y = 91 else
"111111111111" when X = 91 AND Y = 91 else
"111111111111" when X = 92 AND Y = 91 else
"111111111111" when X = 93 AND Y = 91 else
"111111111111" when X = 94 AND Y = 91 else
"111111111111" when X = 95 AND Y = 91 else
"111111111111" when X = 96 AND Y = 91 else
"111111111111" when X = 97 AND Y = 91 else
"111111111111" when X = 98 AND Y = 91 else
"111111111111" when X = 99 AND Y = 91 else
"111111111111" when X = 100 AND Y = 91 else
"111111111111" when X = 101 AND Y = 91 else
"111111111111" when X = 102 AND Y = 91 else
"111111111111" when X = 103 AND Y = 91 else
"111111111111" when X = 104 AND Y = 91 else
"111111111111" when X = 105 AND Y = 91 else
"111111111111" when X = 106 AND Y = 91 else
"111111111111" when X = 107 AND Y = 91 else
"111111111111" when X = 108 AND Y = 91 else
"111111111111" when X = 109 AND Y = 91 else
"111111111111" when X = 110 AND Y = 91 else
"111111111111" when X = 111 AND Y = 91 else
"111111111111" when X = 112 AND Y = 91 else
"111111111111" when X = 113 AND Y = 91 else
"111111111111" when X = 114 AND Y = 91 else
"111111111111" when X = 115 AND Y = 91 else
"111111111111" when X = 116 AND Y = 91 else
"111111111111" when X = 117 AND Y = 91 else
"111111111111" when X = 118 AND Y = 91 else
"111111111111" when X = 119 AND Y = 91 else
"111111111111" when X = 120 AND Y = 91 else
"111111111111" when X = 121 AND Y = 91 else
"111111111111" when X = 122 AND Y = 91 else
"111111111111" when X = 123 AND Y = 91 else
"111111111111" when X = 124 AND Y = 91 else
"111111111111" when X = 125 AND Y = 91 else
"111111111111" when X = 126 AND Y = 91 else
"111111111111" when X = 127 AND Y = 91 else
"111111111111" when X = 128 AND Y = 91 else
"111111111111" when X = 129 AND Y = 91 else
"111111111111" when X = 130 AND Y = 91 else
"111111111111" when X = 131 AND Y = 91 else
"111111111111" when X = 132 AND Y = 91 else
"111111111111" when X = 133 AND Y = 91 else
"111111111111" when X = 134 AND Y = 91 else
"111111111111" when X = 135 AND Y = 91 else
"111111111111" when X = 136 AND Y = 91 else
"111111111111" when X = 137 AND Y = 91 else
"111111111111" when X = 138 AND Y = 91 else
"111111111111" when X = 139 AND Y = 91 else
"111111111111" when X = 140 AND Y = 91 else
"111111111111" when X = 141 AND Y = 91 else
"111111111111" when X = 142 AND Y = 91 else
"111111111111" when X = 143 AND Y = 91 else
"111111111111" when X = 144 AND Y = 91 else
"111111111111" when X = 145 AND Y = 91 else
"111111111111" when X = 146 AND Y = 91 else
"111111111111" when X = 147 AND Y = 91 else
"111111111111" when X = 148 AND Y = 91 else
"111111111111" when X = 149 AND Y = 91 else
"111111111111" when X = 150 AND Y = 91 else
"111111111111" when X = 151 AND Y = 91 else
"111111111111" when X = 152 AND Y = 91 else
"111111111111" when X = 153 AND Y = 91 else
"111111111111" when X = 154 AND Y = 91 else
"111111111111" when X = 155 AND Y = 91 else
"111111111111" when X = 156 AND Y = 91 else
"111111111111" when X = 157 AND Y = 91 else
"111111111111" when X = 158 AND Y = 91 else
"111111111111" when X = 159 AND Y = 91 else
"111111111111" when X = 160 AND Y = 91 else
"111111111111" when X = 161 AND Y = 91 else
"111111111111" when X = 162 AND Y = 91 else
"111111111111" when X = 163 AND Y = 91 else
"111111111111" when X = 164 AND Y = 91 else
"111111111111" when X = 165 AND Y = 91 else
"111111111111" when X = 166 AND Y = 91 else
"111111111111" when X = 167 AND Y = 91 else
"111111111111" when X = 168 AND Y = 91 else
"111111111111" when X = 169 AND Y = 91 else
"111111111111" when X = 170 AND Y = 91 else
"111111111111" when X = 171 AND Y = 91 else
"111111111111" when X = 172 AND Y = 91 else
"111111111111" when X = 173 AND Y = 91 else
"111111111111" when X = 174 AND Y = 91 else
"111111111111" when X = 175 AND Y = 91 else
"111111111111" when X = 176 AND Y = 91 else
"111111111111" when X = 177 AND Y = 91 else
"111111111111" when X = 178 AND Y = 91 else
"111111111111" when X = 179 AND Y = 91 else
"111111111111" when X = 180 AND Y = 91 else
"111111111111" when X = 181 AND Y = 91 else
"111111111111" when X = 182 AND Y = 91 else
"111111111111" when X = 183 AND Y = 91 else
"111111111111" when X = 184 AND Y = 91 else
"111111111111" when X = 185 AND Y = 91 else
"111111111111" when X = 186 AND Y = 91 else
"111111111111" when X = 187 AND Y = 91 else
"111111111111" when X = 188 AND Y = 91 else
"111111111111" when X = 189 AND Y = 91 else
"111111111111" when X = 190 AND Y = 91 else
"111111111111" when X = 191 AND Y = 91 else
"111111111111" when X = 192 AND Y = 91 else
"111111111111" when X = 193 AND Y = 91 else
"111111111111" when X = 194 AND Y = 91 else
"111111111111" when X = 195 AND Y = 91 else
"111111111111" when X = 196 AND Y = 91 else
"111111111111" when X = 197 AND Y = 91 else
"111111111111" when X = 198 AND Y = 91 else
"111111111111" when X = 199 AND Y = 91 else
"111111111111" when X = 200 AND Y = 91 else
"111111111111" when X = 201 AND Y = 91 else
"111111111111" when X = 202 AND Y = 91 else
"111111111111" when X = 203 AND Y = 91 else
"111111111111" when X = 204 AND Y = 91 else
"111111111111" when X = 205 AND Y = 91 else
"111111111111" when X = 206 AND Y = 91 else
"111111111111" when X = 207 AND Y = 91 else
"111111111111" when X = 208 AND Y = 91 else
"111111111111" when X = 209 AND Y = 91 else
"111111111111" when X = 210 AND Y = 91 else
"111111111111" when X = 211 AND Y = 91 else
"111111111111" when X = 212 AND Y = 91 else
"111111111111" when X = 213 AND Y = 91 else
"111111111111" when X = 214 AND Y = 91 else
"111111111111" when X = 215 AND Y = 91 else
"111111111111" when X = 216 AND Y = 91 else
"111111111111" when X = 217 AND Y = 91 else
"111111111111" when X = 218 AND Y = 91 else
"111111111111" when X = 219 AND Y = 91 else
"110111011111" when X = 220 AND Y = 91 else
"110111011111" when X = 221 AND Y = 91 else
"110111011111" when X = 222 AND Y = 91 else
"110111011111" when X = 223 AND Y = 91 else
"110111011111" when X = 224 AND Y = 91 else
"110111011111" when X = 225 AND Y = 91 else
"110111011111" when X = 226 AND Y = 91 else
"110111011111" when X = 227 AND Y = 91 else
"110111011111" when X = 228 AND Y = 91 else
"110111011111" when X = 229 AND Y = 91 else
"111111111111" when X = 230 AND Y = 91 else
"111111111111" when X = 231 AND Y = 91 else
"111111111111" when X = 232 AND Y = 91 else
"111111111111" when X = 233 AND Y = 91 else
"111111111111" when X = 234 AND Y = 91 else
"111111111111" when X = 235 AND Y = 91 else
"111111111111" when X = 236 AND Y = 91 else
"111111111111" when X = 237 AND Y = 91 else
"111111111111" when X = 238 AND Y = 91 else
"111111111111" when X = 239 AND Y = 91 else
"111111111111" when X = 240 AND Y = 91 else
"111111111111" when X = 241 AND Y = 91 else
"111111111111" when X = 242 AND Y = 91 else
"111111111111" when X = 243 AND Y = 91 else
"111111111111" when X = 244 AND Y = 91 else
"111111111111" when X = 245 AND Y = 91 else
"111111111111" when X = 246 AND Y = 91 else
"111111111111" when X = 247 AND Y = 91 else
"111111111111" when X = 248 AND Y = 91 else
"111111111111" when X = 249 AND Y = 91 else
"111111111111" when X = 250 AND Y = 91 else
"111111111111" when X = 251 AND Y = 91 else
"111111111111" when X = 252 AND Y = 91 else
"111111111111" when X = 253 AND Y = 91 else
"111111111111" when X = 254 AND Y = 91 else
"111111111111" when X = 255 AND Y = 91 else
"111111111111" when X = 256 AND Y = 91 else
"111111111111" when X = 257 AND Y = 91 else
"111111111111" when X = 258 AND Y = 91 else
"111111111111" when X = 259 AND Y = 91 else
"111111111111" when X = 260 AND Y = 91 else
"111111111111" when X = 261 AND Y = 91 else
"111111111111" when X = 262 AND Y = 91 else
"111111111111" when X = 263 AND Y = 91 else
"111111111111" when X = 264 AND Y = 91 else
"111111111111" when X = 265 AND Y = 91 else
"111111111111" when X = 266 AND Y = 91 else
"111111111111" when X = 267 AND Y = 91 else
"111111111111" when X = 268 AND Y = 91 else
"111111111111" when X = 269 AND Y = 91 else
"111111111111" when X = 270 AND Y = 91 else
"111111111111" when X = 271 AND Y = 91 else
"111111111111" when X = 272 AND Y = 91 else
"111111111111" when X = 273 AND Y = 91 else
"111111111111" when X = 274 AND Y = 91 else
"110111011111" when X = 275 AND Y = 91 else
"110111011111" when X = 276 AND Y = 91 else
"110111011111" when X = 277 AND Y = 91 else
"110111011111" when X = 278 AND Y = 91 else
"110111011111" when X = 279 AND Y = 91 else
"110111011111" when X = 280 AND Y = 91 else
"110111011111" when X = 281 AND Y = 91 else
"110111011111" when X = 282 AND Y = 91 else
"110111011111" when X = 283 AND Y = 91 else
"110111011111" when X = 284 AND Y = 91 else
"110111011111" when X = 285 AND Y = 91 else
"110111011111" when X = 286 AND Y = 91 else
"110111011111" when X = 287 AND Y = 91 else
"110111011111" when X = 288 AND Y = 91 else
"110111011111" when X = 289 AND Y = 91 else
"110111011111" when X = 290 AND Y = 91 else
"110111011111" when X = 291 AND Y = 91 else
"110111011111" when X = 292 AND Y = 91 else
"110111011111" when X = 293 AND Y = 91 else
"110111011111" when X = 294 AND Y = 91 else
"110111011111" when X = 295 AND Y = 91 else
"110111011111" when X = 296 AND Y = 91 else
"110111011111" when X = 297 AND Y = 91 else
"110111011111" when X = 298 AND Y = 91 else
"110111011111" when X = 299 AND Y = 91 else
"110111011111" when X = 300 AND Y = 91 else
"110111011111" when X = 301 AND Y = 91 else
"110111011111" when X = 302 AND Y = 91 else
"110111011111" when X = 303 AND Y = 91 else
"110111011111" when X = 304 AND Y = 91 else
"110111011111" when X = 305 AND Y = 91 else
"110111011111" when X = 306 AND Y = 91 else
"110111011111" when X = 307 AND Y = 91 else
"110111011111" when X = 308 AND Y = 91 else
"110111011111" when X = 309 AND Y = 91 else
"110111011111" when X = 310 AND Y = 91 else
"110111011111" when X = 311 AND Y = 91 else
"110111011111" when X = 312 AND Y = 91 else
"110111011111" when X = 313 AND Y = 91 else
"110111011111" when X = 314 AND Y = 91 else
"110111011111" when X = 315 AND Y = 91 else
"110111011111" when X = 316 AND Y = 91 else
"110111011111" when X = 317 AND Y = 91 else
"110111011111" when X = 318 AND Y = 91 else
"110111011111" when X = 319 AND Y = 91 else
"000000000000" when X = 320 AND Y = 91 else
"000000000000" when X = 321 AND Y = 91 else
"000000000000" when X = 322 AND Y = 91 else
"000000000000" when X = 323 AND Y = 91 else
"000000000000" when X = 324 AND Y = 91 else
"100010011101" when X = 0 AND Y = 92 else
"100010011101" when X = 1 AND Y = 92 else
"100010011101" when X = 2 AND Y = 92 else
"100010011101" when X = 3 AND Y = 92 else
"100010011101" when X = 4 AND Y = 92 else
"100010011101" when X = 5 AND Y = 92 else
"100010011101" when X = 6 AND Y = 92 else
"100010011101" when X = 7 AND Y = 92 else
"100010011101" when X = 8 AND Y = 92 else
"100010011101" when X = 9 AND Y = 92 else
"100010011101" when X = 10 AND Y = 92 else
"100010011101" when X = 11 AND Y = 92 else
"100010011101" when X = 12 AND Y = 92 else
"100010011101" when X = 13 AND Y = 92 else
"100010011101" when X = 14 AND Y = 92 else
"100010011101" when X = 15 AND Y = 92 else
"100010011101" when X = 16 AND Y = 92 else
"100010011101" when X = 17 AND Y = 92 else
"100010011101" when X = 18 AND Y = 92 else
"100010011101" when X = 19 AND Y = 92 else
"110111011111" when X = 20 AND Y = 92 else
"110111011111" when X = 21 AND Y = 92 else
"110111011111" when X = 22 AND Y = 92 else
"110111011111" when X = 23 AND Y = 92 else
"110111011111" when X = 24 AND Y = 92 else
"110111011111" when X = 25 AND Y = 92 else
"110111011111" when X = 26 AND Y = 92 else
"110111011111" when X = 27 AND Y = 92 else
"110111011111" when X = 28 AND Y = 92 else
"110111011111" when X = 29 AND Y = 92 else
"110111011111" when X = 30 AND Y = 92 else
"110111011111" when X = 31 AND Y = 92 else
"110111011111" when X = 32 AND Y = 92 else
"110111011111" when X = 33 AND Y = 92 else
"110111011111" when X = 34 AND Y = 92 else
"110111011111" when X = 35 AND Y = 92 else
"110111011111" when X = 36 AND Y = 92 else
"110111011111" when X = 37 AND Y = 92 else
"110111011111" when X = 38 AND Y = 92 else
"110111011111" when X = 39 AND Y = 92 else
"110111011111" when X = 40 AND Y = 92 else
"110111011111" when X = 41 AND Y = 92 else
"110111011111" when X = 42 AND Y = 92 else
"110111011111" when X = 43 AND Y = 92 else
"110111011111" when X = 44 AND Y = 92 else
"110111011111" when X = 45 AND Y = 92 else
"110111011111" when X = 46 AND Y = 92 else
"110111011111" when X = 47 AND Y = 92 else
"110111011111" when X = 48 AND Y = 92 else
"110111011111" when X = 49 AND Y = 92 else
"110111011111" when X = 50 AND Y = 92 else
"110111011111" when X = 51 AND Y = 92 else
"110111011111" when X = 52 AND Y = 92 else
"110111011111" when X = 53 AND Y = 92 else
"110111011111" when X = 54 AND Y = 92 else
"110111011111" when X = 55 AND Y = 92 else
"110111011111" when X = 56 AND Y = 92 else
"110111011111" when X = 57 AND Y = 92 else
"110111011111" when X = 58 AND Y = 92 else
"110111011111" when X = 59 AND Y = 92 else
"110111011111" when X = 60 AND Y = 92 else
"110111011111" when X = 61 AND Y = 92 else
"110111011111" when X = 62 AND Y = 92 else
"110111011111" when X = 63 AND Y = 92 else
"110111011111" when X = 64 AND Y = 92 else
"110111011111" when X = 65 AND Y = 92 else
"110111011111" when X = 66 AND Y = 92 else
"110111011111" when X = 67 AND Y = 92 else
"110111011111" when X = 68 AND Y = 92 else
"110111011111" when X = 69 AND Y = 92 else
"111111111111" when X = 70 AND Y = 92 else
"111111111111" when X = 71 AND Y = 92 else
"111111111111" when X = 72 AND Y = 92 else
"111111111111" when X = 73 AND Y = 92 else
"111111111111" when X = 74 AND Y = 92 else
"111111111111" when X = 75 AND Y = 92 else
"111111111111" when X = 76 AND Y = 92 else
"111111111111" when X = 77 AND Y = 92 else
"111111111111" when X = 78 AND Y = 92 else
"111111111111" when X = 79 AND Y = 92 else
"111111111111" when X = 80 AND Y = 92 else
"111111111111" when X = 81 AND Y = 92 else
"111111111111" when X = 82 AND Y = 92 else
"111111111111" when X = 83 AND Y = 92 else
"111111111111" when X = 84 AND Y = 92 else
"111111111111" when X = 85 AND Y = 92 else
"111111111111" when X = 86 AND Y = 92 else
"111111111111" when X = 87 AND Y = 92 else
"111111111111" when X = 88 AND Y = 92 else
"111111111111" when X = 89 AND Y = 92 else
"111111111111" when X = 90 AND Y = 92 else
"111111111111" when X = 91 AND Y = 92 else
"111111111111" when X = 92 AND Y = 92 else
"111111111111" when X = 93 AND Y = 92 else
"111111111111" when X = 94 AND Y = 92 else
"111111111111" when X = 95 AND Y = 92 else
"111111111111" when X = 96 AND Y = 92 else
"111111111111" when X = 97 AND Y = 92 else
"111111111111" when X = 98 AND Y = 92 else
"111111111111" when X = 99 AND Y = 92 else
"111111111111" when X = 100 AND Y = 92 else
"111111111111" when X = 101 AND Y = 92 else
"111111111111" when X = 102 AND Y = 92 else
"111111111111" when X = 103 AND Y = 92 else
"111111111111" when X = 104 AND Y = 92 else
"111111111111" when X = 105 AND Y = 92 else
"111111111111" when X = 106 AND Y = 92 else
"111111111111" when X = 107 AND Y = 92 else
"111111111111" when X = 108 AND Y = 92 else
"111111111111" when X = 109 AND Y = 92 else
"111111111111" when X = 110 AND Y = 92 else
"111111111111" when X = 111 AND Y = 92 else
"111111111111" when X = 112 AND Y = 92 else
"111111111111" when X = 113 AND Y = 92 else
"111111111111" when X = 114 AND Y = 92 else
"111111111111" when X = 115 AND Y = 92 else
"111111111111" when X = 116 AND Y = 92 else
"111111111111" when X = 117 AND Y = 92 else
"111111111111" when X = 118 AND Y = 92 else
"111111111111" when X = 119 AND Y = 92 else
"111111111111" when X = 120 AND Y = 92 else
"111111111111" when X = 121 AND Y = 92 else
"111111111111" when X = 122 AND Y = 92 else
"111111111111" when X = 123 AND Y = 92 else
"111111111111" when X = 124 AND Y = 92 else
"111111111111" when X = 125 AND Y = 92 else
"111111111111" when X = 126 AND Y = 92 else
"111111111111" when X = 127 AND Y = 92 else
"111111111111" when X = 128 AND Y = 92 else
"111111111111" when X = 129 AND Y = 92 else
"111111111111" when X = 130 AND Y = 92 else
"111111111111" when X = 131 AND Y = 92 else
"111111111111" when X = 132 AND Y = 92 else
"111111111111" when X = 133 AND Y = 92 else
"111111111111" when X = 134 AND Y = 92 else
"111111111111" when X = 135 AND Y = 92 else
"111111111111" when X = 136 AND Y = 92 else
"111111111111" when X = 137 AND Y = 92 else
"111111111111" when X = 138 AND Y = 92 else
"111111111111" when X = 139 AND Y = 92 else
"111111111111" when X = 140 AND Y = 92 else
"111111111111" when X = 141 AND Y = 92 else
"111111111111" when X = 142 AND Y = 92 else
"111111111111" when X = 143 AND Y = 92 else
"111111111111" when X = 144 AND Y = 92 else
"111111111111" when X = 145 AND Y = 92 else
"111111111111" when X = 146 AND Y = 92 else
"111111111111" when X = 147 AND Y = 92 else
"111111111111" when X = 148 AND Y = 92 else
"111111111111" when X = 149 AND Y = 92 else
"111111111111" when X = 150 AND Y = 92 else
"111111111111" when X = 151 AND Y = 92 else
"111111111111" when X = 152 AND Y = 92 else
"111111111111" when X = 153 AND Y = 92 else
"111111111111" when X = 154 AND Y = 92 else
"111111111111" when X = 155 AND Y = 92 else
"111111111111" when X = 156 AND Y = 92 else
"111111111111" when X = 157 AND Y = 92 else
"111111111111" when X = 158 AND Y = 92 else
"111111111111" when X = 159 AND Y = 92 else
"111111111111" when X = 160 AND Y = 92 else
"111111111111" when X = 161 AND Y = 92 else
"111111111111" when X = 162 AND Y = 92 else
"111111111111" when X = 163 AND Y = 92 else
"111111111111" when X = 164 AND Y = 92 else
"111111111111" when X = 165 AND Y = 92 else
"111111111111" when X = 166 AND Y = 92 else
"111111111111" when X = 167 AND Y = 92 else
"111111111111" when X = 168 AND Y = 92 else
"111111111111" when X = 169 AND Y = 92 else
"111111111111" when X = 170 AND Y = 92 else
"111111111111" when X = 171 AND Y = 92 else
"111111111111" when X = 172 AND Y = 92 else
"111111111111" when X = 173 AND Y = 92 else
"111111111111" when X = 174 AND Y = 92 else
"111111111111" when X = 175 AND Y = 92 else
"111111111111" when X = 176 AND Y = 92 else
"111111111111" when X = 177 AND Y = 92 else
"111111111111" when X = 178 AND Y = 92 else
"111111111111" when X = 179 AND Y = 92 else
"111111111111" when X = 180 AND Y = 92 else
"111111111111" when X = 181 AND Y = 92 else
"111111111111" when X = 182 AND Y = 92 else
"111111111111" when X = 183 AND Y = 92 else
"111111111111" when X = 184 AND Y = 92 else
"111111111111" when X = 185 AND Y = 92 else
"111111111111" when X = 186 AND Y = 92 else
"111111111111" when X = 187 AND Y = 92 else
"111111111111" when X = 188 AND Y = 92 else
"111111111111" when X = 189 AND Y = 92 else
"111111111111" when X = 190 AND Y = 92 else
"111111111111" when X = 191 AND Y = 92 else
"111111111111" when X = 192 AND Y = 92 else
"111111111111" when X = 193 AND Y = 92 else
"111111111111" when X = 194 AND Y = 92 else
"111111111111" when X = 195 AND Y = 92 else
"111111111111" when X = 196 AND Y = 92 else
"111111111111" when X = 197 AND Y = 92 else
"111111111111" when X = 198 AND Y = 92 else
"111111111111" when X = 199 AND Y = 92 else
"111111111111" when X = 200 AND Y = 92 else
"111111111111" when X = 201 AND Y = 92 else
"111111111111" when X = 202 AND Y = 92 else
"111111111111" when X = 203 AND Y = 92 else
"111111111111" when X = 204 AND Y = 92 else
"111111111111" when X = 205 AND Y = 92 else
"111111111111" when X = 206 AND Y = 92 else
"111111111111" when X = 207 AND Y = 92 else
"111111111111" when X = 208 AND Y = 92 else
"111111111111" when X = 209 AND Y = 92 else
"111111111111" when X = 210 AND Y = 92 else
"111111111111" when X = 211 AND Y = 92 else
"111111111111" when X = 212 AND Y = 92 else
"111111111111" when X = 213 AND Y = 92 else
"111111111111" when X = 214 AND Y = 92 else
"111111111111" when X = 215 AND Y = 92 else
"111111111111" when X = 216 AND Y = 92 else
"111111111111" when X = 217 AND Y = 92 else
"111111111111" when X = 218 AND Y = 92 else
"111111111111" when X = 219 AND Y = 92 else
"110111011111" when X = 220 AND Y = 92 else
"110111011111" when X = 221 AND Y = 92 else
"110111011111" when X = 222 AND Y = 92 else
"110111011111" when X = 223 AND Y = 92 else
"110111011111" when X = 224 AND Y = 92 else
"110111011111" when X = 225 AND Y = 92 else
"110111011111" when X = 226 AND Y = 92 else
"110111011111" when X = 227 AND Y = 92 else
"110111011111" when X = 228 AND Y = 92 else
"110111011111" when X = 229 AND Y = 92 else
"111111111111" when X = 230 AND Y = 92 else
"111111111111" when X = 231 AND Y = 92 else
"111111111111" when X = 232 AND Y = 92 else
"111111111111" when X = 233 AND Y = 92 else
"111111111111" when X = 234 AND Y = 92 else
"111111111111" when X = 235 AND Y = 92 else
"111111111111" when X = 236 AND Y = 92 else
"111111111111" when X = 237 AND Y = 92 else
"111111111111" when X = 238 AND Y = 92 else
"111111111111" when X = 239 AND Y = 92 else
"111111111111" when X = 240 AND Y = 92 else
"111111111111" when X = 241 AND Y = 92 else
"111111111111" when X = 242 AND Y = 92 else
"111111111111" when X = 243 AND Y = 92 else
"111111111111" when X = 244 AND Y = 92 else
"111111111111" when X = 245 AND Y = 92 else
"111111111111" when X = 246 AND Y = 92 else
"111111111111" when X = 247 AND Y = 92 else
"111111111111" when X = 248 AND Y = 92 else
"111111111111" when X = 249 AND Y = 92 else
"111111111111" when X = 250 AND Y = 92 else
"111111111111" when X = 251 AND Y = 92 else
"111111111111" when X = 252 AND Y = 92 else
"111111111111" when X = 253 AND Y = 92 else
"111111111111" when X = 254 AND Y = 92 else
"111111111111" when X = 255 AND Y = 92 else
"111111111111" when X = 256 AND Y = 92 else
"111111111111" when X = 257 AND Y = 92 else
"111111111111" when X = 258 AND Y = 92 else
"111111111111" when X = 259 AND Y = 92 else
"111111111111" when X = 260 AND Y = 92 else
"111111111111" when X = 261 AND Y = 92 else
"111111111111" when X = 262 AND Y = 92 else
"111111111111" when X = 263 AND Y = 92 else
"111111111111" when X = 264 AND Y = 92 else
"111111111111" when X = 265 AND Y = 92 else
"111111111111" when X = 266 AND Y = 92 else
"111111111111" when X = 267 AND Y = 92 else
"111111111111" when X = 268 AND Y = 92 else
"111111111111" when X = 269 AND Y = 92 else
"111111111111" when X = 270 AND Y = 92 else
"111111111111" when X = 271 AND Y = 92 else
"111111111111" when X = 272 AND Y = 92 else
"111111111111" when X = 273 AND Y = 92 else
"111111111111" when X = 274 AND Y = 92 else
"110111011111" when X = 275 AND Y = 92 else
"110111011111" when X = 276 AND Y = 92 else
"110111011111" when X = 277 AND Y = 92 else
"110111011111" when X = 278 AND Y = 92 else
"110111011111" when X = 279 AND Y = 92 else
"110111011111" when X = 280 AND Y = 92 else
"110111011111" when X = 281 AND Y = 92 else
"110111011111" when X = 282 AND Y = 92 else
"110111011111" when X = 283 AND Y = 92 else
"110111011111" when X = 284 AND Y = 92 else
"110111011111" when X = 285 AND Y = 92 else
"110111011111" when X = 286 AND Y = 92 else
"110111011111" when X = 287 AND Y = 92 else
"110111011111" when X = 288 AND Y = 92 else
"110111011111" when X = 289 AND Y = 92 else
"110111011111" when X = 290 AND Y = 92 else
"110111011111" when X = 291 AND Y = 92 else
"110111011111" when X = 292 AND Y = 92 else
"110111011111" when X = 293 AND Y = 92 else
"110111011111" when X = 294 AND Y = 92 else
"110111011111" when X = 295 AND Y = 92 else
"110111011111" when X = 296 AND Y = 92 else
"110111011111" when X = 297 AND Y = 92 else
"110111011111" when X = 298 AND Y = 92 else
"110111011111" when X = 299 AND Y = 92 else
"110111011111" when X = 300 AND Y = 92 else
"110111011111" when X = 301 AND Y = 92 else
"110111011111" when X = 302 AND Y = 92 else
"110111011111" when X = 303 AND Y = 92 else
"110111011111" when X = 304 AND Y = 92 else
"110111011111" when X = 305 AND Y = 92 else
"110111011111" when X = 306 AND Y = 92 else
"110111011111" when X = 307 AND Y = 92 else
"110111011111" when X = 308 AND Y = 92 else
"110111011111" when X = 309 AND Y = 92 else
"110111011111" when X = 310 AND Y = 92 else
"110111011111" when X = 311 AND Y = 92 else
"110111011111" when X = 312 AND Y = 92 else
"110111011111" when X = 313 AND Y = 92 else
"110111011111" when X = 314 AND Y = 92 else
"110111011111" when X = 315 AND Y = 92 else
"110111011111" when X = 316 AND Y = 92 else
"110111011111" when X = 317 AND Y = 92 else
"110111011111" when X = 318 AND Y = 92 else
"110111011111" when X = 319 AND Y = 92 else
"000000000000" when X = 320 AND Y = 92 else
"000000000000" when X = 321 AND Y = 92 else
"000000000000" when X = 322 AND Y = 92 else
"000000000000" when X = 323 AND Y = 92 else
"000000000000" when X = 324 AND Y = 92 else
"100010011101" when X = 0 AND Y = 93 else
"100010011101" when X = 1 AND Y = 93 else
"100010011101" when X = 2 AND Y = 93 else
"100010011101" when X = 3 AND Y = 93 else
"100010011101" when X = 4 AND Y = 93 else
"100010011101" when X = 5 AND Y = 93 else
"100010011101" when X = 6 AND Y = 93 else
"100010011101" when X = 7 AND Y = 93 else
"100010011101" when X = 8 AND Y = 93 else
"100010011101" when X = 9 AND Y = 93 else
"100010011101" when X = 10 AND Y = 93 else
"100010011101" when X = 11 AND Y = 93 else
"100010011101" when X = 12 AND Y = 93 else
"100010011101" when X = 13 AND Y = 93 else
"100010011101" when X = 14 AND Y = 93 else
"100010011101" when X = 15 AND Y = 93 else
"100010011101" when X = 16 AND Y = 93 else
"100010011101" when X = 17 AND Y = 93 else
"100010011101" when X = 18 AND Y = 93 else
"100010011101" when X = 19 AND Y = 93 else
"110111011111" when X = 20 AND Y = 93 else
"110111011111" when X = 21 AND Y = 93 else
"110111011111" when X = 22 AND Y = 93 else
"110111011111" when X = 23 AND Y = 93 else
"110111011111" when X = 24 AND Y = 93 else
"110111011111" when X = 25 AND Y = 93 else
"110111011111" when X = 26 AND Y = 93 else
"110111011111" when X = 27 AND Y = 93 else
"110111011111" when X = 28 AND Y = 93 else
"110111011111" when X = 29 AND Y = 93 else
"110111011111" when X = 30 AND Y = 93 else
"110111011111" when X = 31 AND Y = 93 else
"110111011111" when X = 32 AND Y = 93 else
"110111011111" when X = 33 AND Y = 93 else
"110111011111" when X = 34 AND Y = 93 else
"110111011111" when X = 35 AND Y = 93 else
"110111011111" when X = 36 AND Y = 93 else
"110111011111" when X = 37 AND Y = 93 else
"110111011111" when X = 38 AND Y = 93 else
"110111011111" when X = 39 AND Y = 93 else
"110111011111" when X = 40 AND Y = 93 else
"110111011111" when X = 41 AND Y = 93 else
"110111011111" when X = 42 AND Y = 93 else
"110111011111" when X = 43 AND Y = 93 else
"110111011111" when X = 44 AND Y = 93 else
"110111011111" when X = 45 AND Y = 93 else
"110111011111" when X = 46 AND Y = 93 else
"110111011111" when X = 47 AND Y = 93 else
"110111011111" when X = 48 AND Y = 93 else
"110111011111" when X = 49 AND Y = 93 else
"110111011111" when X = 50 AND Y = 93 else
"110111011111" when X = 51 AND Y = 93 else
"110111011111" when X = 52 AND Y = 93 else
"110111011111" when X = 53 AND Y = 93 else
"110111011111" when X = 54 AND Y = 93 else
"110111011111" when X = 55 AND Y = 93 else
"110111011111" when X = 56 AND Y = 93 else
"110111011111" when X = 57 AND Y = 93 else
"110111011111" when X = 58 AND Y = 93 else
"110111011111" when X = 59 AND Y = 93 else
"110111011111" when X = 60 AND Y = 93 else
"110111011111" when X = 61 AND Y = 93 else
"110111011111" when X = 62 AND Y = 93 else
"110111011111" when X = 63 AND Y = 93 else
"110111011111" when X = 64 AND Y = 93 else
"110111011111" when X = 65 AND Y = 93 else
"110111011111" when X = 66 AND Y = 93 else
"110111011111" when X = 67 AND Y = 93 else
"110111011111" when X = 68 AND Y = 93 else
"110111011111" when X = 69 AND Y = 93 else
"111111111111" when X = 70 AND Y = 93 else
"111111111111" when X = 71 AND Y = 93 else
"111111111111" when X = 72 AND Y = 93 else
"111111111111" when X = 73 AND Y = 93 else
"111111111111" when X = 74 AND Y = 93 else
"111111111111" when X = 75 AND Y = 93 else
"111111111111" when X = 76 AND Y = 93 else
"111111111111" when X = 77 AND Y = 93 else
"111111111111" when X = 78 AND Y = 93 else
"111111111111" when X = 79 AND Y = 93 else
"111111111111" when X = 80 AND Y = 93 else
"111111111111" when X = 81 AND Y = 93 else
"111111111111" when X = 82 AND Y = 93 else
"111111111111" when X = 83 AND Y = 93 else
"111111111111" when X = 84 AND Y = 93 else
"111111111111" when X = 85 AND Y = 93 else
"111111111111" when X = 86 AND Y = 93 else
"111111111111" when X = 87 AND Y = 93 else
"111111111111" when X = 88 AND Y = 93 else
"111111111111" when X = 89 AND Y = 93 else
"111111111111" when X = 90 AND Y = 93 else
"111111111111" when X = 91 AND Y = 93 else
"111111111111" when X = 92 AND Y = 93 else
"111111111111" when X = 93 AND Y = 93 else
"111111111111" when X = 94 AND Y = 93 else
"111111111111" when X = 95 AND Y = 93 else
"111111111111" when X = 96 AND Y = 93 else
"111111111111" when X = 97 AND Y = 93 else
"111111111111" when X = 98 AND Y = 93 else
"111111111111" when X = 99 AND Y = 93 else
"111111111111" when X = 100 AND Y = 93 else
"111111111111" when X = 101 AND Y = 93 else
"111111111111" when X = 102 AND Y = 93 else
"111111111111" when X = 103 AND Y = 93 else
"111111111111" when X = 104 AND Y = 93 else
"111111111111" when X = 105 AND Y = 93 else
"111111111111" when X = 106 AND Y = 93 else
"111111111111" when X = 107 AND Y = 93 else
"111111111111" when X = 108 AND Y = 93 else
"111111111111" when X = 109 AND Y = 93 else
"111111111111" when X = 110 AND Y = 93 else
"111111111111" when X = 111 AND Y = 93 else
"111111111111" when X = 112 AND Y = 93 else
"111111111111" when X = 113 AND Y = 93 else
"111111111111" when X = 114 AND Y = 93 else
"111111111111" when X = 115 AND Y = 93 else
"111111111111" when X = 116 AND Y = 93 else
"111111111111" when X = 117 AND Y = 93 else
"111111111111" when X = 118 AND Y = 93 else
"111111111111" when X = 119 AND Y = 93 else
"111111111111" when X = 120 AND Y = 93 else
"111111111111" when X = 121 AND Y = 93 else
"111111111111" when X = 122 AND Y = 93 else
"111111111111" when X = 123 AND Y = 93 else
"111111111111" when X = 124 AND Y = 93 else
"111111111111" when X = 125 AND Y = 93 else
"111111111111" when X = 126 AND Y = 93 else
"111111111111" when X = 127 AND Y = 93 else
"111111111111" when X = 128 AND Y = 93 else
"111111111111" when X = 129 AND Y = 93 else
"111111111111" when X = 130 AND Y = 93 else
"111111111111" when X = 131 AND Y = 93 else
"111111111111" when X = 132 AND Y = 93 else
"111111111111" when X = 133 AND Y = 93 else
"111111111111" when X = 134 AND Y = 93 else
"111111111111" when X = 135 AND Y = 93 else
"111111111111" when X = 136 AND Y = 93 else
"111111111111" when X = 137 AND Y = 93 else
"111111111111" when X = 138 AND Y = 93 else
"111111111111" when X = 139 AND Y = 93 else
"111111111111" when X = 140 AND Y = 93 else
"111111111111" when X = 141 AND Y = 93 else
"111111111111" when X = 142 AND Y = 93 else
"111111111111" when X = 143 AND Y = 93 else
"111111111111" when X = 144 AND Y = 93 else
"111111111111" when X = 145 AND Y = 93 else
"111111111111" when X = 146 AND Y = 93 else
"111111111111" when X = 147 AND Y = 93 else
"111111111111" when X = 148 AND Y = 93 else
"111111111111" when X = 149 AND Y = 93 else
"111111111111" when X = 150 AND Y = 93 else
"111111111111" when X = 151 AND Y = 93 else
"111111111111" when X = 152 AND Y = 93 else
"111111111111" when X = 153 AND Y = 93 else
"111111111111" when X = 154 AND Y = 93 else
"111111111111" when X = 155 AND Y = 93 else
"111111111111" when X = 156 AND Y = 93 else
"111111111111" when X = 157 AND Y = 93 else
"111111111111" when X = 158 AND Y = 93 else
"111111111111" when X = 159 AND Y = 93 else
"111111111111" when X = 160 AND Y = 93 else
"111111111111" when X = 161 AND Y = 93 else
"111111111111" when X = 162 AND Y = 93 else
"111111111111" when X = 163 AND Y = 93 else
"111111111111" when X = 164 AND Y = 93 else
"111111111111" when X = 165 AND Y = 93 else
"111111111111" when X = 166 AND Y = 93 else
"111111111111" when X = 167 AND Y = 93 else
"111111111111" when X = 168 AND Y = 93 else
"111111111111" when X = 169 AND Y = 93 else
"111111111111" when X = 170 AND Y = 93 else
"111111111111" when X = 171 AND Y = 93 else
"111111111111" when X = 172 AND Y = 93 else
"111111111111" when X = 173 AND Y = 93 else
"111111111111" when X = 174 AND Y = 93 else
"111111111111" when X = 175 AND Y = 93 else
"111111111111" when X = 176 AND Y = 93 else
"111111111111" when X = 177 AND Y = 93 else
"111111111111" when X = 178 AND Y = 93 else
"111111111111" when X = 179 AND Y = 93 else
"111111111111" when X = 180 AND Y = 93 else
"111111111111" when X = 181 AND Y = 93 else
"111111111111" when X = 182 AND Y = 93 else
"111111111111" when X = 183 AND Y = 93 else
"111111111111" when X = 184 AND Y = 93 else
"111111111111" when X = 185 AND Y = 93 else
"111111111111" when X = 186 AND Y = 93 else
"111111111111" when X = 187 AND Y = 93 else
"111111111111" when X = 188 AND Y = 93 else
"111111111111" when X = 189 AND Y = 93 else
"111111111111" when X = 190 AND Y = 93 else
"111111111111" when X = 191 AND Y = 93 else
"111111111111" when X = 192 AND Y = 93 else
"111111111111" when X = 193 AND Y = 93 else
"111111111111" when X = 194 AND Y = 93 else
"111111111111" when X = 195 AND Y = 93 else
"111111111111" when X = 196 AND Y = 93 else
"111111111111" when X = 197 AND Y = 93 else
"111111111111" when X = 198 AND Y = 93 else
"111111111111" when X = 199 AND Y = 93 else
"111111111111" when X = 200 AND Y = 93 else
"111111111111" when X = 201 AND Y = 93 else
"111111111111" when X = 202 AND Y = 93 else
"111111111111" when X = 203 AND Y = 93 else
"111111111111" when X = 204 AND Y = 93 else
"111111111111" when X = 205 AND Y = 93 else
"111111111111" when X = 206 AND Y = 93 else
"111111111111" when X = 207 AND Y = 93 else
"111111111111" when X = 208 AND Y = 93 else
"111111111111" when X = 209 AND Y = 93 else
"111111111111" when X = 210 AND Y = 93 else
"111111111111" when X = 211 AND Y = 93 else
"111111111111" when X = 212 AND Y = 93 else
"111111111111" when X = 213 AND Y = 93 else
"111111111111" when X = 214 AND Y = 93 else
"111111111111" when X = 215 AND Y = 93 else
"111111111111" when X = 216 AND Y = 93 else
"111111111111" when X = 217 AND Y = 93 else
"111111111111" when X = 218 AND Y = 93 else
"111111111111" when X = 219 AND Y = 93 else
"110111011111" when X = 220 AND Y = 93 else
"110111011111" when X = 221 AND Y = 93 else
"110111011111" when X = 222 AND Y = 93 else
"110111011111" when X = 223 AND Y = 93 else
"110111011111" when X = 224 AND Y = 93 else
"110111011111" when X = 225 AND Y = 93 else
"110111011111" when X = 226 AND Y = 93 else
"110111011111" when X = 227 AND Y = 93 else
"110111011111" when X = 228 AND Y = 93 else
"110111011111" when X = 229 AND Y = 93 else
"111111111111" when X = 230 AND Y = 93 else
"111111111111" when X = 231 AND Y = 93 else
"111111111111" when X = 232 AND Y = 93 else
"111111111111" when X = 233 AND Y = 93 else
"111111111111" when X = 234 AND Y = 93 else
"111111111111" when X = 235 AND Y = 93 else
"111111111111" when X = 236 AND Y = 93 else
"111111111111" when X = 237 AND Y = 93 else
"111111111111" when X = 238 AND Y = 93 else
"111111111111" when X = 239 AND Y = 93 else
"111111111111" when X = 240 AND Y = 93 else
"111111111111" when X = 241 AND Y = 93 else
"111111111111" when X = 242 AND Y = 93 else
"111111111111" when X = 243 AND Y = 93 else
"111111111111" when X = 244 AND Y = 93 else
"111111111111" when X = 245 AND Y = 93 else
"111111111111" when X = 246 AND Y = 93 else
"111111111111" when X = 247 AND Y = 93 else
"111111111111" when X = 248 AND Y = 93 else
"111111111111" when X = 249 AND Y = 93 else
"111111111111" when X = 250 AND Y = 93 else
"111111111111" when X = 251 AND Y = 93 else
"111111111111" when X = 252 AND Y = 93 else
"111111111111" when X = 253 AND Y = 93 else
"111111111111" when X = 254 AND Y = 93 else
"111111111111" when X = 255 AND Y = 93 else
"111111111111" when X = 256 AND Y = 93 else
"111111111111" when X = 257 AND Y = 93 else
"111111111111" when X = 258 AND Y = 93 else
"111111111111" when X = 259 AND Y = 93 else
"111111111111" when X = 260 AND Y = 93 else
"111111111111" when X = 261 AND Y = 93 else
"111111111111" when X = 262 AND Y = 93 else
"111111111111" when X = 263 AND Y = 93 else
"111111111111" when X = 264 AND Y = 93 else
"111111111111" when X = 265 AND Y = 93 else
"111111111111" when X = 266 AND Y = 93 else
"111111111111" when X = 267 AND Y = 93 else
"111111111111" when X = 268 AND Y = 93 else
"111111111111" when X = 269 AND Y = 93 else
"111111111111" when X = 270 AND Y = 93 else
"111111111111" when X = 271 AND Y = 93 else
"111111111111" when X = 272 AND Y = 93 else
"111111111111" when X = 273 AND Y = 93 else
"111111111111" when X = 274 AND Y = 93 else
"110111011111" when X = 275 AND Y = 93 else
"110111011111" when X = 276 AND Y = 93 else
"110111011111" when X = 277 AND Y = 93 else
"110111011111" when X = 278 AND Y = 93 else
"110111011111" when X = 279 AND Y = 93 else
"110111011111" when X = 280 AND Y = 93 else
"110111011111" when X = 281 AND Y = 93 else
"110111011111" when X = 282 AND Y = 93 else
"110111011111" when X = 283 AND Y = 93 else
"110111011111" when X = 284 AND Y = 93 else
"110111011111" when X = 285 AND Y = 93 else
"110111011111" when X = 286 AND Y = 93 else
"110111011111" when X = 287 AND Y = 93 else
"110111011111" when X = 288 AND Y = 93 else
"110111011111" when X = 289 AND Y = 93 else
"110111011111" when X = 290 AND Y = 93 else
"110111011111" when X = 291 AND Y = 93 else
"110111011111" when X = 292 AND Y = 93 else
"110111011111" when X = 293 AND Y = 93 else
"110111011111" when X = 294 AND Y = 93 else
"110111011111" when X = 295 AND Y = 93 else
"110111011111" when X = 296 AND Y = 93 else
"110111011111" when X = 297 AND Y = 93 else
"110111011111" when X = 298 AND Y = 93 else
"110111011111" when X = 299 AND Y = 93 else
"110111011111" when X = 300 AND Y = 93 else
"110111011111" when X = 301 AND Y = 93 else
"110111011111" when X = 302 AND Y = 93 else
"110111011111" when X = 303 AND Y = 93 else
"110111011111" when X = 304 AND Y = 93 else
"110111011111" when X = 305 AND Y = 93 else
"110111011111" when X = 306 AND Y = 93 else
"110111011111" when X = 307 AND Y = 93 else
"110111011111" when X = 308 AND Y = 93 else
"110111011111" when X = 309 AND Y = 93 else
"110111011111" when X = 310 AND Y = 93 else
"110111011111" when X = 311 AND Y = 93 else
"110111011111" when X = 312 AND Y = 93 else
"110111011111" when X = 313 AND Y = 93 else
"110111011111" when X = 314 AND Y = 93 else
"110111011111" when X = 315 AND Y = 93 else
"110111011111" when X = 316 AND Y = 93 else
"110111011111" when X = 317 AND Y = 93 else
"110111011111" when X = 318 AND Y = 93 else
"110111011111" when X = 319 AND Y = 93 else
"000000000000" when X = 320 AND Y = 93 else
"000000000000" when X = 321 AND Y = 93 else
"000000000000" when X = 322 AND Y = 93 else
"000000000000" when X = 323 AND Y = 93 else
"000000000000" when X = 324 AND Y = 93 else
"100010011101" when X = 0 AND Y = 94 else
"100010011101" when X = 1 AND Y = 94 else
"100010011101" when X = 2 AND Y = 94 else
"100010011101" when X = 3 AND Y = 94 else
"100010011101" when X = 4 AND Y = 94 else
"100010011101" when X = 5 AND Y = 94 else
"100010011101" when X = 6 AND Y = 94 else
"100010011101" when X = 7 AND Y = 94 else
"100010011101" when X = 8 AND Y = 94 else
"100010011101" when X = 9 AND Y = 94 else
"100010011101" when X = 10 AND Y = 94 else
"100010011101" when X = 11 AND Y = 94 else
"100010011101" when X = 12 AND Y = 94 else
"100010011101" when X = 13 AND Y = 94 else
"100010011101" when X = 14 AND Y = 94 else
"100010011101" when X = 15 AND Y = 94 else
"100010011101" when X = 16 AND Y = 94 else
"100010011101" when X = 17 AND Y = 94 else
"100010011101" when X = 18 AND Y = 94 else
"100010011101" when X = 19 AND Y = 94 else
"110111011111" when X = 20 AND Y = 94 else
"110111011111" when X = 21 AND Y = 94 else
"110111011111" when X = 22 AND Y = 94 else
"110111011111" when X = 23 AND Y = 94 else
"110111011111" when X = 24 AND Y = 94 else
"110111011111" when X = 25 AND Y = 94 else
"110111011111" when X = 26 AND Y = 94 else
"110111011111" when X = 27 AND Y = 94 else
"110111011111" when X = 28 AND Y = 94 else
"110111011111" when X = 29 AND Y = 94 else
"110111011111" when X = 30 AND Y = 94 else
"110111011111" when X = 31 AND Y = 94 else
"110111011111" when X = 32 AND Y = 94 else
"110111011111" when X = 33 AND Y = 94 else
"110111011111" when X = 34 AND Y = 94 else
"110111011111" when X = 35 AND Y = 94 else
"110111011111" when X = 36 AND Y = 94 else
"110111011111" when X = 37 AND Y = 94 else
"110111011111" when X = 38 AND Y = 94 else
"110111011111" when X = 39 AND Y = 94 else
"110111011111" when X = 40 AND Y = 94 else
"110111011111" when X = 41 AND Y = 94 else
"110111011111" when X = 42 AND Y = 94 else
"110111011111" when X = 43 AND Y = 94 else
"110111011111" when X = 44 AND Y = 94 else
"110111011111" when X = 45 AND Y = 94 else
"110111011111" when X = 46 AND Y = 94 else
"110111011111" when X = 47 AND Y = 94 else
"110111011111" when X = 48 AND Y = 94 else
"110111011111" when X = 49 AND Y = 94 else
"110111011111" when X = 50 AND Y = 94 else
"110111011111" when X = 51 AND Y = 94 else
"110111011111" when X = 52 AND Y = 94 else
"110111011111" when X = 53 AND Y = 94 else
"110111011111" when X = 54 AND Y = 94 else
"110111011111" when X = 55 AND Y = 94 else
"110111011111" when X = 56 AND Y = 94 else
"110111011111" when X = 57 AND Y = 94 else
"110111011111" when X = 58 AND Y = 94 else
"110111011111" when X = 59 AND Y = 94 else
"110111011111" when X = 60 AND Y = 94 else
"110111011111" when X = 61 AND Y = 94 else
"110111011111" when X = 62 AND Y = 94 else
"110111011111" when X = 63 AND Y = 94 else
"110111011111" when X = 64 AND Y = 94 else
"110111011111" when X = 65 AND Y = 94 else
"110111011111" when X = 66 AND Y = 94 else
"110111011111" when X = 67 AND Y = 94 else
"110111011111" when X = 68 AND Y = 94 else
"110111011111" when X = 69 AND Y = 94 else
"111111111111" when X = 70 AND Y = 94 else
"111111111111" when X = 71 AND Y = 94 else
"111111111111" when X = 72 AND Y = 94 else
"111111111111" when X = 73 AND Y = 94 else
"111111111111" when X = 74 AND Y = 94 else
"111111111111" when X = 75 AND Y = 94 else
"111111111111" when X = 76 AND Y = 94 else
"111111111111" when X = 77 AND Y = 94 else
"111111111111" when X = 78 AND Y = 94 else
"111111111111" when X = 79 AND Y = 94 else
"111111111111" when X = 80 AND Y = 94 else
"111111111111" when X = 81 AND Y = 94 else
"111111111111" when X = 82 AND Y = 94 else
"111111111111" when X = 83 AND Y = 94 else
"111111111111" when X = 84 AND Y = 94 else
"111111111111" when X = 85 AND Y = 94 else
"111111111111" when X = 86 AND Y = 94 else
"111111111111" when X = 87 AND Y = 94 else
"111111111111" when X = 88 AND Y = 94 else
"111111111111" when X = 89 AND Y = 94 else
"111111111111" when X = 90 AND Y = 94 else
"111111111111" when X = 91 AND Y = 94 else
"111111111111" when X = 92 AND Y = 94 else
"111111111111" when X = 93 AND Y = 94 else
"111111111111" when X = 94 AND Y = 94 else
"111111111111" when X = 95 AND Y = 94 else
"111111111111" when X = 96 AND Y = 94 else
"111111111111" when X = 97 AND Y = 94 else
"111111111111" when X = 98 AND Y = 94 else
"111111111111" when X = 99 AND Y = 94 else
"111111111111" when X = 100 AND Y = 94 else
"111111111111" when X = 101 AND Y = 94 else
"111111111111" when X = 102 AND Y = 94 else
"111111111111" when X = 103 AND Y = 94 else
"111111111111" when X = 104 AND Y = 94 else
"111111111111" when X = 105 AND Y = 94 else
"111111111111" when X = 106 AND Y = 94 else
"111111111111" when X = 107 AND Y = 94 else
"111111111111" when X = 108 AND Y = 94 else
"111111111111" when X = 109 AND Y = 94 else
"111111111111" when X = 110 AND Y = 94 else
"111111111111" when X = 111 AND Y = 94 else
"111111111111" when X = 112 AND Y = 94 else
"111111111111" when X = 113 AND Y = 94 else
"111111111111" when X = 114 AND Y = 94 else
"111111111111" when X = 115 AND Y = 94 else
"111111111111" when X = 116 AND Y = 94 else
"111111111111" when X = 117 AND Y = 94 else
"111111111111" when X = 118 AND Y = 94 else
"111111111111" when X = 119 AND Y = 94 else
"111111111111" when X = 120 AND Y = 94 else
"111111111111" when X = 121 AND Y = 94 else
"111111111111" when X = 122 AND Y = 94 else
"111111111111" when X = 123 AND Y = 94 else
"111111111111" when X = 124 AND Y = 94 else
"111111111111" when X = 125 AND Y = 94 else
"111111111111" when X = 126 AND Y = 94 else
"111111111111" when X = 127 AND Y = 94 else
"111111111111" when X = 128 AND Y = 94 else
"111111111111" when X = 129 AND Y = 94 else
"111111111111" when X = 130 AND Y = 94 else
"111111111111" when X = 131 AND Y = 94 else
"111111111111" when X = 132 AND Y = 94 else
"111111111111" when X = 133 AND Y = 94 else
"111111111111" when X = 134 AND Y = 94 else
"111111111111" when X = 135 AND Y = 94 else
"111111111111" when X = 136 AND Y = 94 else
"111111111111" when X = 137 AND Y = 94 else
"111111111111" when X = 138 AND Y = 94 else
"111111111111" when X = 139 AND Y = 94 else
"111111111111" when X = 140 AND Y = 94 else
"111111111111" when X = 141 AND Y = 94 else
"111111111111" when X = 142 AND Y = 94 else
"111111111111" when X = 143 AND Y = 94 else
"111111111111" when X = 144 AND Y = 94 else
"111111111111" when X = 145 AND Y = 94 else
"111111111111" when X = 146 AND Y = 94 else
"111111111111" when X = 147 AND Y = 94 else
"111111111111" when X = 148 AND Y = 94 else
"111111111111" when X = 149 AND Y = 94 else
"111111111111" when X = 150 AND Y = 94 else
"111111111111" when X = 151 AND Y = 94 else
"111111111111" when X = 152 AND Y = 94 else
"111111111111" when X = 153 AND Y = 94 else
"111111111111" when X = 154 AND Y = 94 else
"111111111111" when X = 155 AND Y = 94 else
"111111111111" when X = 156 AND Y = 94 else
"111111111111" when X = 157 AND Y = 94 else
"111111111111" when X = 158 AND Y = 94 else
"111111111111" when X = 159 AND Y = 94 else
"111111111111" when X = 160 AND Y = 94 else
"111111111111" when X = 161 AND Y = 94 else
"111111111111" when X = 162 AND Y = 94 else
"111111111111" when X = 163 AND Y = 94 else
"111111111111" when X = 164 AND Y = 94 else
"111111111111" when X = 165 AND Y = 94 else
"111111111111" when X = 166 AND Y = 94 else
"111111111111" when X = 167 AND Y = 94 else
"111111111111" when X = 168 AND Y = 94 else
"111111111111" when X = 169 AND Y = 94 else
"111111111111" when X = 170 AND Y = 94 else
"111111111111" when X = 171 AND Y = 94 else
"111111111111" when X = 172 AND Y = 94 else
"111111111111" when X = 173 AND Y = 94 else
"111111111111" when X = 174 AND Y = 94 else
"111111111111" when X = 175 AND Y = 94 else
"111111111111" when X = 176 AND Y = 94 else
"111111111111" when X = 177 AND Y = 94 else
"111111111111" when X = 178 AND Y = 94 else
"111111111111" when X = 179 AND Y = 94 else
"111111111111" when X = 180 AND Y = 94 else
"111111111111" when X = 181 AND Y = 94 else
"111111111111" when X = 182 AND Y = 94 else
"111111111111" when X = 183 AND Y = 94 else
"111111111111" when X = 184 AND Y = 94 else
"111111111111" when X = 185 AND Y = 94 else
"111111111111" when X = 186 AND Y = 94 else
"111111111111" when X = 187 AND Y = 94 else
"111111111111" when X = 188 AND Y = 94 else
"111111111111" when X = 189 AND Y = 94 else
"111111111111" when X = 190 AND Y = 94 else
"111111111111" when X = 191 AND Y = 94 else
"111111111111" when X = 192 AND Y = 94 else
"111111111111" when X = 193 AND Y = 94 else
"111111111111" when X = 194 AND Y = 94 else
"111111111111" when X = 195 AND Y = 94 else
"111111111111" when X = 196 AND Y = 94 else
"111111111111" when X = 197 AND Y = 94 else
"111111111111" when X = 198 AND Y = 94 else
"111111111111" when X = 199 AND Y = 94 else
"111111111111" when X = 200 AND Y = 94 else
"111111111111" when X = 201 AND Y = 94 else
"111111111111" when X = 202 AND Y = 94 else
"111111111111" when X = 203 AND Y = 94 else
"111111111111" when X = 204 AND Y = 94 else
"111111111111" when X = 205 AND Y = 94 else
"111111111111" when X = 206 AND Y = 94 else
"111111111111" when X = 207 AND Y = 94 else
"111111111111" when X = 208 AND Y = 94 else
"111111111111" when X = 209 AND Y = 94 else
"111111111111" when X = 210 AND Y = 94 else
"111111111111" when X = 211 AND Y = 94 else
"111111111111" when X = 212 AND Y = 94 else
"111111111111" when X = 213 AND Y = 94 else
"111111111111" when X = 214 AND Y = 94 else
"111111111111" when X = 215 AND Y = 94 else
"111111111111" when X = 216 AND Y = 94 else
"111111111111" when X = 217 AND Y = 94 else
"111111111111" when X = 218 AND Y = 94 else
"111111111111" when X = 219 AND Y = 94 else
"110111011111" when X = 220 AND Y = 94 else
"110111011111" when X = 221 AND Y = 94 else
"110111011111" when X = 222 AND Y = 94 else
"110111011111" when X = 223 AND Y = 94 else
"110111011111" when X = 224 AND Y = 94 else
"110111011111" when X = 225 AND Y = 94 else
"110111011111" when X = 226 AND Y = 94 else
"110111011111" when X = 227 AND Y = 94 else
"110111011111" when X = 228 AND Y = 94 else
"110111011111" when X = 229 AND Y = 94 else
"111111111111" when X = 230 AND Y = 94 else
"111111111111" when X = 231 AND Y = 94 else
"111111111111" when X = 232 AND Y = 94 else
"111111111111" when X = 233 AND Y = 94 else
"111111111111" when X = 234 AND Y = 94 else
"111111111111" when X = 235 AND Y = 94 else
"111111111111" when X = 236 AND Y = 94 else
"111111111111" when X = 237 AND Y = 94 else
"111111111111" when X = 238 AND Y = 94 else
"111111111111" when X = 239 AND Y = 94 else
"111111111111" when X = 240 AND Y = 94 else
"111111111111" when X = 241 AND Y = 94 else
"111111111111" when X = 242 AND Y = 94 else
"111111111111" when X = 243 AND Y = 94 else
"111111111111" when X = 244 AND Y = 94 else
"111111111111" when X = 245 AND Y = 94 else
"111111111111" when X = 246 AND Y = 94 else
"111111111111" when X = 247 AND Y = 94 else
"111111111111" when X = 248 AND Y = 94 else
"111111111111" when X = 249 AND Y = 94 else
"111111111111" when X = 250 AND Y = 94 else
"111111111111" when X = 251 AND Y = 94 else
"111111111111" when X = 252 AND Y = 94 else
"111111111111" when X = 253 AND Y = 94 else
"111111111111" when X = 254 AND Y = 94 else
"111111111111" when X = 255 AND Y = 94 else
"111111111111" when X = 256 AND Y = 94 else
"111111111111" when X = 257 AND Y = 94 else
"111111111111" when X = 258 AND Y = 94 else
"111111111111" when X = 259 AND Y = 94 else
"111111111111" when X = 260 AND Y = 94 else
"111111111111" when X = 261 AND Y = 94 else
"111111111111" when X = 262 AND Y = 94 else
"111111111111" when X = 263 AND Y = 94 else
"111111111111" when X = 264 AND Y = 94 else
"111111111111" when X = 265 AND Y = 94 else
"111111111111" when X = 266 AND Y = 94 else
"111111111111" when X = 267 AND Y = 94 else
"111111111111" when X = 268 AND Y = 94 else
"111111111111" when X = 269 AND Y = 94 else
"111111111111" when X = 270 AND Y = 94 else
"111111111111" when X = 271 AND Y = 94 else
"111111111111" when X = 272 AND Y = 94 else
"111111111111" when X = 273 AND Y = 94 else
"111111111111" when X = 274 AND Y = 94 else
"110111011111" when X = 275 AND Y = 94 else
"110111011111" when X = 276 AND Y = 94 else
"110111011111" when X = 277 AND Y = 94 else
"110111011111" when X = 278 AND Y = 94 else
"110111011111" when X = 279 AND Y = 94 else
"110111011111" when X = 280 AND Y = 94 else
"110111011111" when X = 281 AND Y = 94 else
"110111011111" when X = 282 AND Y = 94 else
"110111011111" when X = 283 AND Y = 94 else
"110111011111" when X = 284 AND Y = 94 else
"110111011111" when X = 285 AND Y = 94 else
"110111011111" when X = 286 AND Y = 94 else
"110111011111" when X = 287 AND Y = 94 else
"110111011111" when X = 288 AND Y = 94 else
"110111011111" when X = 289 AND Y = 94 else
"110111011111" when X = 290 AND Y = 94 else
"110111011111" when X = 291 AND Y = 94 else
"110111011111" when X = 292 AND Y = 94 else
"110111011111" when X = 293 AND Y = 94 else
"110111011111" when X = 294 AND Y = 94 else
"110111011111" when X = 295 AND Y = 94 else
"110111011111" when X = 296 AND Y = 94 else
"110111011111" when X = 297 AND Y = 94 else
"110111011111" when X = 298 AND Y = 94 else
"110111011111" when X = 299 AND Y = 94 else
"110111011111" when X = 300 AND Y = 94 else
"110111011111" when X = 301 AND Y = 94 else
"110111011111" when X = 302 AND Y = 94 else
"110111011111" when X = 303 AND Y = 94 else
"110111011111" when X = 304 AND Y = 94 else
"110111011111" when X = 305 AND Y = 94 else
"110111011111" when X = 306 AND Y = 94 else
"110111011111" when X = 307 AND Y = 94 else
"110111011111" when X = 308 AND Y = 94 else
"110111011111" when X = 309 AND Y = 94 else
"110111011111" when X = 310 AND Y = 94 else
"110111011111" when X = 311 AND Y = 94 else
"110111011111" when X = 312 AND Y = 94 else
"110111011111" when X = 313 AND Y = 94 else
"110111011111" when X = 314 AND Y = 94 else
"110111011111" when X = 315 AND Y = 94 else
"110111011111" when X = 316 AND Y = 94 else
"110111011111" when X = 317 AND Y = 94 else
"110111011111" when X = 318 AND Y = 94 else
"110111011111" when X = 319 AND Y = 94 else
"000000000000" when X = 320 AND Y = 94 else
"000000000000" when X = 321 AND Y = 94 else
"000000000000" when X = 322 AND Y = 94 else
"000000000000" when X = 323 AND Y = 94 else
"000000000000" when X = 324 AND Y = 94 else
"100010011101" when X = 0 AND Y = 95 else
"100010011101" when X = 1 AND Y = 95 else
"100010011101" when X = 2 AND Y = 95 else
"100010011101" when X = 3 AND Y = 95 else
"100010011101" when X = 4 AND Y = 95 else
"100010011101" when X = 5 AND Y = 95 else
"100010011101" when X = 6 AND Y = 95 else
"100010011101" when X = 7 AND Y = 95 else
"100010011101" when X = 8 AND Y = 95 else
"100010011101" when X = 9 AND Y = 95 else
"100010011101" when X = 10 AND Y = 95 else
"100010011101" when X = 11 AND Y = 95 else
"100010011101" when X = 12 AND Y = 95 else
"100010011101" when X = 13 AND Y = 95 else
"100010011101" when X = 14 AND Y = 95 else
"110111011111" when X = 15 AND Y = 95 else
"110111011111" when X = 16 AND Y = 95 else
"110111011111" when X = 17 AND Y = 95 else
"110111011111" when X = 18 AND Y = 95 else
"110111011111" when X = 19 AND Y = 95 else
"110111011111" when X = 20 AND Y = 95 else
"110111011111" when X = 21 AND Y = 95 else
"110111011111" when X = 22 AND Y = 95 else
"110111011111" when X = 23 AND Y = 95 else
"110111011111" when X = 24 AND Y = 95 else
"110111011111" when X = 25 AND Y = 95 else
"110111011111" when X = 26 AND Y = 95 else
"110111011111" when X = 27 AND Y = 95 else
"110111011111" when X = 28 AND Y = 95 else
"110111011111" when X = 29 AND Y = 95 else
"110111011111" when X = 30 AND Y = 95 else
"110111011111" when X = 31 AND Y = 95 else
"110111011111" when X = 32 AND Y = 95 else
"110111011111" when X = 33 AND Y = 95 else
"110111011111" when X = 34 AND Y = 95 else
"110111011111" when X = 35 AND Y = 95 else
"110111011111" when X = 36 AND Y = 95 else
"110111011111" when X = 37 AND Y = 95 else
"110111011111" when X = 38 AND Y = 95 else
"110111011111" when X = 39 AND Y = 95 else
"110111011111" when X = 40 AND Y = 95 else
"110111011111" when X = 41 AND Y = 95 else
"110111011111" when X = 42 AND Y = 95 else
"110111011111" when X = 43 AND Y = 95 else
"110111011111" when X = 44 AND Y = 95 else
"110111011111" when X = 45 AND Y = 95 else
"110111011111" when X = 46 AND Y = 95 else
"110111011111" when X = 47 AND Y = 95 else
"110111011111" when X = 48 AND Y = 95 else
"110111011111" when X = 49 AND Y = 95 else
"110111011111" when X = 50 AND Y = 95 else
"110111011111" when X = 51 AND Y = 95 else
"110111011111" when X = 52 AND Y = 95 else
"110111011111" when X = 53 AND Y = 95 else
"110111011111" when X = 54 AND Y = 95 else
"110111011111" when X = 55 AND Y = 95 else
"110111011111" when X = 56 AND Y = 95 else
"110111011111" when X = 57 AND Y = 95 else
"110111011111" when X = 58 AND Y = 95 else
"110111011111" when X = 59 AND Y = 95 else
"110111011111" when X = 60 AND Y = 95 else
"110111011111" when X = 61 AND Y = 95 else
"110111011111" when X = 62 AND Y = 95 else
"110111011111" when X = 63 AND Y = 95 else
"110111011111" when X = 64 AND Y = 95 else
"110111011111" when X = 65 AND Y = 95 else
"110111011111" when X = 66 AND Y = 95 else
"110111011111" when X = 67 AND Y = 95 else
"110111011111" when X = 68 AND Y = 95 else
"110111011111" when X = 69 AND Y = 95 else
"111111111111" when X = 70 AND Y = 95 else
"111111111111" when X = 71 AND Y = 95 else
"111111111111" when X = 72 AND Y = 95 else
"111111111111" when X = 73 AND Y = 95 else
"111111111111" when X = 74 AND Y = 95 else
"111111111111" when X = 75 AND Y = 95 else
"111111111111" when X = 76 AND Y = 95 else
"111111111111" when X = 77 AND Y = 95 else
"111111111111" when X = 78 AND Y = 95 else
"111111111111" when X = 79 AND Y = 95 else
"111111111111" when X = 80 AND Y = 95 else
"111111111111" when X = 81 AND Y = 95 else
"111111111111" when X = 82 AND Y = 95 else
"111111111111" when X = 83 AND Y = 95 else
"111111111111" when X = 84 AND Y = 95 else
"111111111111" when X = 85 AND Y = 95 else
"111111111111" when X = 86 AND Y = 95 else
"111111111111" when X = 87 AND Y = 95 else
"111111111111" when X = 88 AND Y = 95 else
"111111111111" when X = 89 AND Y = 95 else
"111111111111" when X = 90 AND Y = 95 else
"111111111111" when X = 91 AND Y = 95 else
"111111111111" when X = 92 AND Y = 95 else
"111111111111" when X = 93 AND Y = 95 else
"111111111111" when X = 94 AND Y = 95 else
"111111111111" when X = 95 AND Y = 95 else
"111111111111" when X = 96 AND Y = 95 else
"111111111111" when X = 97 AND Y = 95 else
"111111111111" when X = 98 AND Y = 95 else
"111111111111" when X = 99 AND Y = 95 else
"111111111111" when X = 100 AND Y = 95 else
"111111111111" when X = 101 AND Y = 95 else
"111111111111" when X = 102 AND Y = 95 else
"111111111111" when X = 103 AND Y = 95 else
"111111111111" when X = 104 AND Y = 95 else
"111111111111" when X = 105 AND Y = 95 else
"111111111111" when X = 106 AND Y = 95 else
"111111111111" when X = 107 AND Y = 95 else
"111111111111" when X = 108 AND Y = 95 else
"111111111111" when X = 109 AND Y = 95 else
"111111111111" when X = 110 AND Y = 95 else
"111111111111" when X = 111 AND Y = 95 else
"111111111111" when X = 112 AND Y = 95 else
"111111111111" when X = 113 AND Y = 95 else
"111111111111" when X = 114 AND Y = 95 else
"111111111111" when X = 115 AND Y = 95 else
"111111111111" when X = 116 AND Y = 95 else
"111111111111" when X = 117 AND Y = 95 else
"111111111111" when X = 118 AND Y = 95 else
"111111111111" when X = 119 AND Y = 95 else
"111111111111" when X = 120 AND Y = 95 else
"111111111111" when X = 121 AND Y = 95 else
"111111111111" when X = 122 AND Y = 95 else
"111111111111" when X = 123 AND Y = 95 else
"111111111111" when X = 124 AND Y = 95 else
"111111111111" when X = 125 AND Y = 95 else
"111111111111" when X = 126 AND Y = 95 else
"111111111111" when X = 127 AND Y = 95 else
"111111111111" when X = 128 AND Y = 95 else
"111111111111" when X = 129 AND Y = 95 else
"111111111111" when X = 130 AND Y = 95 else
"111111111111" when X = 131 AND Y = 95 else
"111111111111" when X = 132 AND Y = 95 else
"111111111111" when X = 133 AND Y = 95 else
"111111111111" when X = 134 AND Y = 95 else
"111111111111" when X = 135 AND Y = 95 else
"111111111111" when X = 136 AND Y = 95 else
"111111111111" when X = 137 AND Y = 95 else
"111111111111" when X = 138 AND Y = 95 else
"111111111111" when X = 139 AND Y = 95 else
"111111111111" when X = 140 AND Y = 95 else
"111111111111" when X = 141 AND Y = 95 else
"111111111111" when X = 142 AND Y = 95 else
"111111111111" when X = 143 AND Y = 95 else
"111111111111" when X = 144 AND Y = 95 else
"111111111111" when X = 145 AND Y = 95 else
"111111111111" when X = 146 AND Y = 95 else
"111111111111" when X = 147 AND Y = 95 else
"111111111111" when X = 148 AND Y = 95 else
"111111111111" when X = 149 AND Y = 95 else
"111111111111" when X = 150 AND Y = 95 else
"111111111111" when X = 151 AND Y = 95 else
"111111111111" when X = 152 AND Y = 95 else
"111111111111" when X = 153 AND Y = 95 else
"111111111111" when X = 154 AND Y = 95 else
"111111111111" when X = 155 AND Y = 95 else
"111111111111" when X = 156 AND Y = 95 else
"111111111111" when X = 157 AND Y = 95 else
"111111111111" when X = 158 AND Y = 95 else
"111111111111" when X = 159 AND Y = 95 else
"111111111111" when X = 160 AND Y = 95 else
"111111111111" when X = 161 AND Y = 95 else
"111111111111" when X = 162 AND Y = 95 else
"111111111111" when X = 163 AND Y = 95 else
"111111111111" when X = 164 AND Y = 95 else
"111111111111" when X = 165 AND Y = 95 else
"111111111111" when X = 166 AND Y = 95 else
"111111111111" when X = 167 AND Y = 95 else
"111111111111" when X = 168 AND Y = 95 else
"111111111111" when X = 169 AND Y = 95 else
"111111111111" when X = 170 AND Y = 95 else
"111111111111" when X = 171 AND Y = 95 else
"111111111111" when X = 172 AND Y = 95 else
"111111111111" when X = 173 AND Y = 95 else
"111111111111" when X = 174 AND Y = 95 else
"111111111111" when X = 175 AND Y = 95 else
"111111111111" when X = 176 AND Y = 95 else
"111111111111" when X = 177 AND Y = 95 else
"111111111111" when X = 178 AND Y = 95 else
"111111111111" when X = 179 AND Y = 95 else
"111111111111" when X = 180 AND Y = 95 else
"111111111111" when X = 181 AND Y = 95 else
"111111111111" when X = 182 AND Y = 95 else
"111111111111" when X = 183 AND Y = 95 else
"111111111111" when X = 184 AND Y = 95 else
"111111111111" when X = 185 AND Y = 95 else
"111111111111" when X = 186 AND Y = 95 else
"111111111111" when X = 187 AND Y = 95 else
"111111111111" when X = 188 AND Y = 95 else
"111111111111" when X = 189 AND Y = 95 else
"111111111111" when X = 190 AND Y = 95 else
"111111111111" when X = 191 AND Y = 95 else
"111111111111" when X = 192 AND Y = 95 else
"111111111111" when X = 193 AND Y = 95 else
"111111111111" when X = 194 AND Y = 95 else
"111111111111" when X = 195 AND Y = 95 else
"111111111111" when X = 196 AND Y = 95 else
"111111111111" when X = 197 AND Y = 95 else
"111111111111" when X = 198 AND Y = 95 else
"111111111111" when X = 199 AND Y = 95 else
"111111111111" when X = 200 AND Y = 95 else
"111111111111" when X = 201 AND Y = 95 else
"111111111111" when X = 202 AND Y = 95 else
"111111111111" when X = 203 AND Y = 95 else
"111111111111" when X = 204 AND Y = 95 else
"110111011111" when X = 205 AND Y = 95 else
"110111011111" when X = 206 AND Y = 95 else
"110111011111" when X = 207 AND Y = 95 else
"110111011111" when X = 208 AND Y = 95 else
"110111011111" when X = 209 AND Y = 95 else
"110111011111" when X = 210 AND Y = 95 else
"110111011111" when X = 211 AND Y = 95 else
"110111011111" when X = 212 AND Y = 95 else
"110111011111" when X = 213 AND Y = 95 else
"110111011111" when X = 214 AND Y = 95 else
"110111011111" when X = 215 AND Y = 95 else
"110111011111" when X = 216 AND Y = 95 else
"110111011111" when X = 217 AND Y = 95 else
"110111011111" when X = 218 AND Y = 95 else
"110111011111" when X = 219 AND Y = 95 else
"111111111111" when X = 220 AND Y = 95 else
"111111111111" when X = 221 AND Y = 95 else
"111111111111" when X = 222 AND Y = 95 else
"111111111111" when X = 223 AND Y = 95 else
"111111111111" when X = 224 AND Y = 95 else
"111111111111" when X = 225 AND Y = 95 else
"111111111111" when X = 226 AND Y = 95 else
"111111111111" when X = 227 AND Y = 95 else
"111111111111" when X = 228 AND Y = 95 else
"111111111111" when X = 229 AND Y = 95 else
"111111111111" when X = 230 AND Y = 95 else
"111111111111" when X = 231 AND Y = 95 else
"111111111111" when X = 232 AND Y = 95 else
"111111111111" when X = 233 AND Y = 95 else
"111111111111" when X = 234 AND Y = 95 else
"111111111111" when X = 235 AND Y = 95 else
"111111111111" when X = 236 AND Y = 95 else
"111111111111" when X = 237 AND Y = 95 else
"111111111111" when X = 238 AND Y = 95 else
"111111111111" when X = 239 AND Y = 95 else
"111111111111" when X = 240 AND Y = 95 else
"111111111111" when X = 241 AND Y = 95 else
"111111111111" when X = 242 AND Y = 95 else
"111111111111" when X = 243 AND Y = 95 else
"111111111111" when X = 244 AND Y = 95 else
"111111111111" when X = 245 AND Y = 95 else
"111111111111" when X = 246 AND Y = 95 else
"111111111111" when X = 247 AND Y = 95 else
"111111111111" when X = 248 AND Y = 95 else
"111111111111" when X = 249 AND Y = 95 else
"111111111111" when X = 250 AND Y = 95 else
"111111111111" when X = 251 AND Y = 95 else
"111111111111" when X = 252 AND Y = 95 else
"111111111111" when X = 253 AND Y = 95 else
"111111111111" when X = 254 AND Y = 95 else
"111111111111" when X = 255 AND Y = 95 else
"111111111111" when X = 256 AND Y = 95 else
"111111111111" when X = 257 AND Y = 95 else
"111111111111" when X = 258 AND Y = 95 else
"111111111111" when X = 259 AND Y = 95 else
"111111111111" when X = 260 AND Y = 95 else
"111111111111" when X = 261 AND Y = 95 else
"111111111111" when X = 262 AND Y = 95 else
"111111111111" when X = 263 AND Y = 95 else
"111111111111" when X = 264 AND Y = 95 else
"111111111111" when X = 265 AND Y = 95 else
"111111111111" when X = 266 AND Y = 95 else
"111111111111" when X = 267 AND Y = 95 else
"111111111111" when X = 268 AND Y = 95 else
"111111111111" when X = 269 AND Y = 95 else
"111111111111" when X = 270 AND Y = 95 else
"111111111111" when X = 271 AND Y = 95 else
"111111111111" when X = 272 AND Y = 95 else
"111111111111" when X = 273 AND Y = 95 else
"111111111111" when X = 274 AND Y = 95 else
"110111011111" when X = 275 AND Y = 95 else
"110111011111" when X = 276 AND Y = 95 else
"110111011111" when X = 277 AND Y = 95 else
"110111011111" when X = 278 AND Y = 95 else
"110111011111" when X = 279 AND Y = 95 else
"110111011111" when X = 280 AND Y = 95 else
"110111011111" when X = 281 AND Y = 95 else
"110111011111" when X = 282 AND Y = 95 else
"110111011111" when X = 283 AND Y = 95 else
"110111011111" when X = 284 AND Y = 95 else
"111111111111" when X = 285 AND Y = 95 else
"111111111111" when X = 286 AND Y = 95 else
"111111111111" when X = 287 AND Y = 95 else
"111111111111" when X = 288 AND Y = 95 else
"111111111111" when X = 289 AND Y = 95 else
"111111111111" when X = 290 AND Y = 95 else
"111111111111" when X = 291 AND Y = 95 else
"111111111111" when X = 292 AND Y = 95 else
"111111111111" when X = 293 AND Y = 95 else
"111111111111" when X = 294 AND Y = 95 else
"111111111111" when X = 295 AND Y = 95 else
"111111111111" when X = 296 AND Y = 95 else
"111111111111" when X = 297 AND Y = 95 else
"111111111111" when X = 298 AND Y = 95 else
"111111111111" when X = 299 AND Y = 95 else
"111111111111" when X = 300 AND Y = 95 else
"111111111111" when X = 301 AND Y = 95 else
"111111111111" when X = 302 AND Y = 95 else
"111111111111" when X = 303 AND Y = 95 else
"111111111111" when X = 304 AND Y = 95 else
"110111011111" when X = 305 AND Y = 95 else
"110111011111" when X = 306 AND Y = 95 else
"110111011111" when X = 307 AND Y = 95 else
"110111011111" when X = 308 AND Y = 95 else
"110111011111" when X = 309 AND Y = 95 else
"110111011111" when X = 310 AND Y = 95 else
"110111011111" when X = 311 AND Y = 95 else
"110111011111" when X = 312 AND Y = 95 else
"110111011111" when X = 313 AND Y = 95 else
"110111011111" when X = 314 AND Y = 95 else
"110111011111" when X = 315 AND Y = 95 else
"110111011111" when X = 316 AND Y = 95 else
"110111011111" when X = 317 AND Y = 95 else
"110111011111" when X = 318 AND Y = 95 else
"110111011111" when X = 319 AND Y = 95 else
"110111011111" when X = 320 AND Y = 95 else
"110111011111" when X = 321 AND Y = 95 else
"110111011111" when X = 322 AND Y = 95 else
"110111011111" when X = 323 AND Y = 95 else
"110111011111" when X = 324 AND Y = 95 else
"100010011101" when X = 0 AND Y = 96 else
"100010011101" when X = 1 AND Y = 96 else
"100010011101" when X = 2 AND Y = 96 else
"100010011101" when X = 3 AND Y = 96 else
"100010011101" when X = 4 AND Y = 96 else
"100010011101" when X = 5 AND Y = 96 else
"100010011101" when X = 6 AND Y = 96 else
"100010011101" when X = 7 AND Y = 96 else
"100010011101" when X = 8 AND Y = 96 else
"100010011101" when X = 9 AND Y = 96 else
"100010011101" when X = 10 AND Y = 96 else
"100010011101" when X = 11 AND Y = 96 else
"100010011101" when X = 12 AND Y = 96 else
"100010011101" when X = 13 AND Y = 96 else
"100010011101" when X = 14 AND Y = 96 else
"110111011111" when X = 15 AND Y = 96 else
"110111011111" when X = 16 AND Y = 96 else
"110111011111" when X = 17 AND Y = 96 else
"110111011111" when X = 18 AND Y = 96 else
"110111011111" when X = 19 AND Y = 96 else
"110111011111" when X = 20 AND Y = 96 else
"110111011111" when X = 21 AND Y = 96 else
"110111011111" when X = 22 AND Y = 96 else
"110111011111" when X = 23 AND Y = 96 else
"110111011111" when X = 24 AND Y = 96 else
"110111011111" when X = 25 AND Y = 96 else
"110111011111" when X = 26 AND Y = 96 else
"110111011111" when X = 27 AND Y = 96 else
"110111011111" when X = 28 AND Y = 96 else
"110111011111" when X = 29 AND Y = 96 else
"110111011111" when X = 30 AND Y = 96 else
"110111011111" when X = 31 AND Y = 96 else
"110111011111" when X = 32 AND Y = 96 else
"110111011111" when X = 33 AND Y = 96 else
"110111011111" when X = 34 AND Y = 96 else
"110111011111" when X = 35 AND Y = 96 else
"110111011111" when X = 36 AND Y = 96 else
"110111011111" when X = 37 AND Y = 96 else
"110111011111" when X = 38 AND Y = 96 else
"110111011111" when X = 39 AND Y = 96 else
"110111011111" when X = 40 AND Y = 96 else
"110111011111" when X = 41 AND Y = 96 else
"110111011111" when X = 42 AND Y = 96 else
"110111011111" when X = 43 AND Y = 96 else
"110111011111" when X = 44 AND Y = 96 else
"110111011111" when X = 45 AND Y = 96 else
"110111011111" when X = 46 AND Y = 96 else
"110111011111" when X = 47 AND Y = 96 else
"110111011111" when X = 48 AND Y = 96 else
"110111011111" when X = 49 AND Y = 96 else
"110111011111" when X = 50 AND Y = 96 else
"110111011111" when X = 51 AND Y = 96 else
"110111011111" when X = 52 AND Y = 96 else
"110111011111" when X = 53 AND Y = 96 else
"110111011111" when X = 54 AND Y = 96 else
"110111011111" when X = 55 AND Y = 96 else
"110111011111" when X = 56 AND Y = 96 else
"110111011111" when X = 57 AND Y = 96 else
"110111011111" when X = 58 AND Y = 96 else
"110111011111" when X = 59 AND Y = 96 else
"110111011111" when X = 60 AND Y = 96 else
"110111011111" when X = 61 AND Y = 96 else
"110111011111" when X = 62 AND Y = 96 else
"110111011111" when X = 63 AND Y = 96 else
"110111011111" when X = 64 AND Y = 96 else
"110111011111" when X = 65 AND Y = 96 else
"110111011111" when X = 66 AND Y = 96 else
"110111011111" when X = 67 AND Y = 96 else
"110111011111" when X = 68 AND Y = 96 else
"110111011111" when X = 69 AND Y = 96 else
"111111111111" when X = 70 AND Y = 96 else
"111111111111" when X = 71 AND Y = 96 else
"111111111111" when X = 72 AND Y = 96 else
"111111111111" when X = 73 AND Y = 96 else
"111111111111" when X = 74 AND Y = 96 else
"111111111111" when X = 75 AND Y = 96 else
"111111111111" when X = 76 AND Y = 96 else
"111111111111" when X = 77 AND Y = 96 else
"111111111111" when X = 78 AND Y = 96 else
"111111111111" when X = 79 AND Y = 96 else
"111111111111" when X = 80 AND Y = 96 else
"111111111111" when X = 81 AND Y = 96 else
"111111111111" when X = 82 AND Y = 96 else
"111111111111" when X = 83 AND Y = 96 else
"111111111111" when X = 84 AND Y = 96 else
"111111111111" when X = 85 AND Y = 96 else
"111111111111" when X = 86 AND Y = 96 else
"111111111111" when X = 87 AND Y = 96 else
"111111111111" when X = 88 AND Y = 96 else
"111111111111" when X = 89 AND Y = 96 else
"111111111111" when X = 90 AND Y = 96 else
"111111111111" when X = 91 AND Y = 96 else
"111111111111" when X = 92 AND Y = 96 else
"111111111111" when X = 93 AND Y = 96 else
"111111111111" when X = 94 AND Y = 96 else
"111111111111" when X = 95 AND Y = 96 else
"111111111111" when X = 96 AND Y = 96 else
"111111111111" when X = 97 AND Y = 96 else
"111111111111" when X = 98 AND Y = 96 else
"111111111111" when X = 99 AND Y = 96 else
"111111111111" when X = 100 AND Y = 96 else
"111111111111" when X = 101 AND Y = 96 else
"111111111111" when X = 102 AND Y = 96 else
"111111111111" when X = 103 AND Y = 96 else
"111111111111" when X = 104 AND Y = 96 else
"111111111111" when X = 105 AND Y = 96 else
"111111111111" when X = 106 AND Y = 96 else
"111111111111" when X = 107 AND Y = 96 else
"111111111111" when X = 108 AND Y = 96 else
"111111111111" when X = 109 AND Y = 96 else
"111111111111" when X = 110 AND Y = 96 else
"111111111111" when X = 111 AND Y = 96 else
"111111111111" when X = 112 AND Y = 96 else
"111111111111" when X = 113 AND Y = 96 else
"111111111111" when X = 114 AND Y = 96 else
"111111111111" when X = 115 AND Y = 96 else
"111111111111" when X = 116 AND Y = 96 else
"111111111111" when X = 117 AND Y = 96 else
"111111111111" when X = 118 AND Y = 96 else
"111111111111" when X = 119 AND Y = 96 else
"111111111111" when X = 120 AND Y = 96 else
"111111111111" when X = 121 AND Y = 96 else
"111111111111" when X = 122 AND Y = 96 else
"111111111111" when X = 123 AND Y = 96 else
"111111111111" when X = 124 AND Y = 96 else
"111111111111" when X = 125 AND Y = 96 else
"111111111111" when X = 126 AND Y = 96 else
"111111111111" when X = 127 AND Y = 96 else
"111111111111" when X = 128 AND Y = 96 else
"111111111111" when X = 129 AND Y = 96 else
"111111111111" when X = 130 AND Y = 96 else
"111111111111" when X = 131 AND Y = 96 else
"111111111111" when X = 132 AND Y = 96 else
"111111111111" when X = 133 AND Y = 96 else
"111111111111" when X = 134 AND Y = 96 else
"111111111111" when X = 135 AND Y = 96 else
"111111111111" when X = 136 AND Y = 96 else
"111111111111" when X = 137 AND Y = 96 else
"111111111111" when X = 138 AND Y = 96 else
"111111111111" when X = 139 AND Y = 96 else
"111111111111" when X = 140 AND Y = 96 else
"111111111111" when X = 141 AND Y = 96 else
"111111111111" when X = 142 AND Y = 96 else
"111111111111" when X = 143 AND Y = 96 else
"111111111111" when X = 144 AND Y = 96 else
"111111111111" when X = 145 AND Y = 96 else
"111111111111" when X = 146 AND Y = 96 else
"111111111111" when X = 147 AND Y = 96 else
"111111111111" when X = 148 AND Y = 96 else
"111111111111" when X = 149 AND Y = 96 else
"111111111111" when X = 150 AND Y = 96 else
"111111111111" when X = 151 AND Y = 96 else
"111111111111" when X = 152 AND Y = 96 else
"111111111111" when X = 153 AND Y = 96 else
"111111111111" when X = 154 AND Y = 96 else
"111111111111" when X = 155 AND Y = 96 else
"111111111111" when X = 156 AND Y = 96 else
"111111111111" when X = 157 AND Y = 96 else
"111111111111" when X = 158 AND Y = 96 else
"111111111111" when X = 159 AND Y = 96 else
"111111111111" when X = 160 AND Y = 96 else
"111111111111" when X = 161 AND Y = 96 else
"111111111111" when X = 162 AND Y = 96 else
"111111111111" when X = 163 AND Y = 96 else
"111111111111" when X = 164 AND Y = 96 else
"111111111111" when X = 165 AND Y = 96 else
"111111111111" when X = 166 AND Y = 96 else
"111111111111" when X = 167 AND Y = 96 else
"111111111111" when X = 168 AND Y = 96 else
"111111111111" when X = 169 AND Y = 96 else
"111111111111" when X = 170 AND Y = 96 else
"111111111111" when X = 171 AND Y = 96 else
"111111111111" when X = 172 AND Y = 96 else
"111111111111" when X = 173 AND Y = 96 else
"111111111111" when X = 174 AND Y = 96 else
"111111111111" when X = 175 AND Y = 96 else
"111111111111" when X = 176 AND Y = 96 else
"111111111111" when X = 177 AND Y = 96 else
"111111111111" when X = 178 AND Y = 96 else
"111111111111" when X = 179 AND Y = 96 else
"111111111111" when X = 180 AND Y = 96 else
"111111111111" when X = 181 AND Y = 96 else
"111111111111" when X = 182 AND Y = 96 else
"111111111111" when X = 183 AND Y = 96 else
"111111111111" when X = 184 AND Y = 96 else
"111111111111" when X = 185 AND Y = 96 else
"111111111111" when X = 186 AND Y = 96 else
"111111111111" when X = 187 AND Y = 96 else
"111111111111" when X = 188 AND Y = 96 else
"111111111111" when X = 189 AND Y = 96 else
"111111111111" when X = 190 AND Y = 96 else
"111111111111" when X = 191 AND Y = 96 else
"111111111111" when X = 192 AND Y = 96 else
"111111111111" when X = 193 AND Y = 96 else
"111111111111" when X = 194 AND Y = 96 else
"111111111111" when X = 195 AND Y = 96 else
"111111111111" when X = 196 AND Y = 96 else
"111111111111" when X = 197 AND Y = 96 else
"111111111111" when X = 198 AND Y = 96 else
"111111111111" when X = 199 AND Y = 96 else
"111111111111" when X = 200 AND Y = 96 else
"111111111111" when X = 201 AND Y = 96 else
"111111111111" when X = 202 AND Y = 96 else
"111111111111" when X = 203 AND Y = 96 else
"111111111111" when X = 204 AND Y = 96 else
"110111011111" when X = 205 AND Y = 96 else
"110111011111" when X = 206 AND Y = 96 else
"110111011111" when X = 207 AND Y = 96 else
"110111011111" when X = 208 AND Y = 96 else
"110111011111" when X = 209 AND Y = 96 else
"110111011111" when X = 210 AND Y = 96 else
"110111011111" when X = 211 AND Y = 96 else
"110111011111" when X = 212 AND Y = 96 else
"110111011111" when X = 213 AND Y = 96 else
"110111011111" when X = 214 AND Y = 96 else
"110111011111" when X = 215 AND Y = 96 else
"110111011111" when X = 216 AND Y = 96 else
"110111011111" when X = 217 AND Y = 96 else
"110111011111" when X = 218 AND Y = 96 else
"110111011111" when X = 219 AND Y = 96 else
"111111111111" when X = 220 AND Y = 96 else
"111111111111" when X = 221 AND Y = 96 else
"111111111111" when X = 222 AND Y = 96 else
"111111111111" when X = 223 AND Y = 96 else
"111111111111" when X = 224 AND Y = 96 else
"111111111111" when X = 225 AND Y = 96 else
"111111111111" when X = 226 AND Y = 96 else
"111111111111" when X = 227 AND Y = 96 else
"111111111111" when X = 228 AND Y = 96 else
"111111111111" when X = 229 AND Y = 96 else
"111111111111" when X = 230 AND Y = 96 else
"111111111111" when X = 231 AND Y = 96 else
"111111111111" when X = 232 AND Y = 96 else
"111111111111" when X = 233 AND Y = 96 else
"111111111111" when X = 234 AND Y = 96 else
"111111111111" when X = 235 AND Y = 96 else
"111111111111" when X = 236 AND Y = 96 else
"111111111111" when X = 237 AND Y = 96 else
"111111111111" when X = 238 AND Y = 96 else
"111111111111" when X = 239 AND Y = 96 else
"111111111111" when X = 240 AND Y = 96 else
"111111111111" when X = 241 AND Y = 96 else
"111111111111" when X = 242 AND Y = 96 else
"111111111111" when X = 243 AND Y = 96 else
"111111111111" when X = 244 AND Y = 96 else
"111111111111" when X = 245 AND Y = 96 else
"111111111111" when X = 246 AND Y = 96 else
"111111111111" when X = 247 AND Y = 96 else
"111111111111" when X = 248 AND Y = 96 else
"111111111111" when X = 249 AND Y = 96 else
"111111111111" when X = 250 AND Y = 96 else
"111111111111" when X = 251 AND Y = 96 else
"111111111111" when X = 252 AND Y = 96 else
"111111111111" when X = 253 AND Y = 96 else
"111111111111" when X = 254 AND Y = 96 else
"111111111111" when X = 255 AND Y = 96 else
"111111111111" when X = 256 AND Y = 96 else
"111111111111" when X = 257 AND Y = 96 else
"111111111111" when X = 258 AND Y = 96 else
"111111111111" when X = 259 AND Y = 96 else
"111111111111" when X = 260 AND Y = 96 else
"111111111111" when X = 261 AND Y = 96 else
"111111111111" when X = 262 AND Y = 96 else
"111111111111" when X = 263 AND Y = 96 else
"111111111111" when X = 264 AND Y = 96 else
"111111111111" when X = 265 AND Y = 96 else
"111111111111" when X = 266 AND Y = 96 else
"111111111111" when X = 267 AND Y = 96 else
"111111111111" when X = 268 AND Y = 96 else
"111111111111" when X = 269 AND Y = 96 else
"111111111111" when X = 270 AND Y = 96 else
"111111111111" when X = 271 AND Y = 96 else
"111111111111" when X = 272 AND Y = 96 else
"111111111111" when X = 273 AND Y = 96 else
"111111111111" when X = 274 AND Y = 96 else
"110111011111" when X = 275 AND Y = 96 else
"110111011111" when X = 276 AND Y = 96 else
"110111011111" when X = 277 AND Y = 96 else
"110111011111" when X = 278 AND Y = 96 else
"110111011111" when X = 279 AND Y = 96 else
"110111011111" when X = 280 AND Y = 96 else
"110111011111" when X = 281 AND Y = 96 else
"110111011111" when X = 282 AND Y = 96 else
"110111011111" when X = 283 AND Y = 96 else
"110111011111" when X = 284 AND Y = 96 else
"111111111111" when X = 285 AND Y = 96 else
"111111111111" when X = 286 AND Y = 96 else
"111111111111" when X = 287 AND Y = 96 else
"111111111111" when X = 288 AND Y = 96 else
"111111111111" when X = 289 AND Y = 96 else
"111111111111" when X = 290 AND Y = 96 else
"111111111111" when X = 291 AND Y = 96 else
"111111111111" when X = 292 AND Y = 96 else
"111111111111" when X = 293 AND Y = 96 else
"111111111111" when X = 294 AND Y = 96 else
"111111111111" when X = 295 AND Y = 96 else
"111111111111" when X = 296 AND Y = 96 else
"111111111111" when X = 297 AND Y = 96 else
"111111111111" when X = 298 AND Y = 96 else
"111111111111" when X = 299 AND Y = 96 else
"111111111111" when X = 300 AND Y = 96 else
"111111111111" when X = 301 AND Y = 96 else
"111111111111" when X = 302 AND Y = 96 else
"111111111111" when X = 303 AND Y = 96 else
"111111111111" when X = 304 AND Y = 96 else
"110111011111" when X = 305 AND Y = 96 else
"110111011111" when X = 306 AND Y = 96 else
"110111011111" when X = 307 AND Y = 96 else
"110111011111" when X = 308 AND Y = 96 else
"110111011111" when X = 309 AND Y = 96 else
"110111011111" when X = 310 AND Y = 96 else
"110111011111" when X = 311 AND Y = 96 else
"110111011111" when X = 312 AND Y = 96 else
"110111011111" when X = 313 AND Y = 96 else
"110111011111" when X = 314 AND Y = 96 else
"110111011111" when X = 315 AND Y = 96 else
"110111011111" when X = 316 AND Y = 96 else
"110111011111" when X = 317 AND Y = 96 else
"110111011111" when X = 318 AND Y = 96 else
"110111011111" when X = 319 AND Y = 96 else
"110111011111" when X = 320 AND Y = 96 else
"110111011111" when X = 321 AND Y = 96 else
"110111011111" when X = 322 AND Y = 96 else
"110111011111" when X = 323 AND Y = 96 else
"110111011111" when X = 324 AND Y = 96 else
"100010011101" when X = 0 AND Y = 97 else
"100010011101" when X = 1 AND Y = 97 else
"100010011101" when X = 2 AND Y = 97 else
"100010011101" when X = 3 AND Y = 97 else
"100010011101" when X = 4 AND Y = 97 else
"100010011101" when X = 5 AND Y = 97 else
"100010011101" when X = 6 AND Y = 97 else
"100010011101" when X = 7 AND Y = 97 else
"100010011101" when X = 8 AND Y = 97 else
"100010011101" when X = 9 AND Y = 97 else
"100010011101" when X = 10 AND Y = 97 else
"100010011101" when X = 11 AND Y = 97 else
"100010011101" when X = 12 AND Y = 97 else
"100010011101" when X = 13 AND Y = 97 else
"100010011101" when X = 14 AND Y = 97 else
"110111011111" when X = 15 AND Y = 97 else
"110111011111" when X = 16 AND Y = 97 else
"110111011111" when X = 17 AND Y = 97 else
"110111011111" when X = 18 AND Y = 97 else
"110111011111" when X = 19 AND Y = 97 else
"110111011111" when X = 20 AND Y = 97 else
"110111011111" when X = 21 AND Y = 97 else
"110111011111" when X = 22 AND Y = 97 else
"110111011111" when X = 23 AND Y = 97 else
"110111011111" when X = 24 AND Y = 97 else
"110111011111" when X = 25 AND Y = 97 else
"110111011111" when X = 26 AND Y = 97 else
"110111011111" when X = 27 AND Y = 97 else
"110111011111" when X = 28 AND Y = 97 else
"110111011111" when X = 29 AND Y = 97 else
"110111011111" when X = 30 AND Y = 97 else
"110111011111" when X = 31 AND Y = 97 else
"110111011111" when X = 32 AND Y = 97 else
"110111011111" when X = 33 AND Y = 97 else
"110111011111" when X = 34 AND Y = 97 else
"110111011111" when X = 35 AND Y = 97 else
"110111011111" when X = 36 AND Y = 97 else
"110111011111" when X = 37 AND Y = 97 else
"110111011111" when X = 38 AND Y = 97 else
"110111011111" when X = 39 AND Y = 97 else
"110111011111" when X = 40 AND Y = 97 else
"110111011111" when X = 41 AND Y = 97 else
"110111011111" when X = 42 AND Y = 97 else
"110111011111" when X = 43 AND Y = 97 else
"110111011111" when X = 44 AND Y = 97 else
"110111011111" when X = 45 AND Y = 97 else
"110111011111" when X = 46 AND Y = 97 else
"110111011111" when X = 47 AND Y = 97 else
"110111011111" when X = 48 AND Y = 97 else
"110111011111" when X = 49 AND Y = 97 else
"110111011111" when X = 50 AND Y = 97 else
"110111011111" when X = 51 AND Y = 97 else
"110111011111" when X = 52 AND Y = 97 else
"110111011111" when X = 53 AND Y = 97 else
"110111011111" when X = 54 AND Y = 97 else
"110111011111" when X = 55 AND Y = 97 else
"110111011111" when X = 56 AND Y = 97 else
"110111011111" when X = 57 AND Y = 97 else
"110111011111" when X = 58 AND Y = 97 else
"110111011111" when X = 59 AND Y = 97 else
"110111011111" when X = 60 AND Y = 97 else
"110111011111" when X = 61 AND Y = 97 else
"110111011111" when X = 62 AND Y = 97 else
"110111011111" when X = 63 AND Y = 97 else
"110111011111" when X = 64 AND Y = 97 else
"110111011111" when X = 65 AND Y = 97 else
"110111011111" when X = 66 AND Y = 97 else
"110111011111" when X = 67 AND Y = 97 else
"110111011111" when X = 68 AND Y = 97 else
"110111011111" when X = 69 AND Y = 97 else
"111111111111" when X = 70 AND Y = 97 else
"111111111111" when X = 71 AND Y = 97 else
"111111111111" when X = 72 AND Y = 97 else
"111111111111" when X = 73 AND Y = 97 else
"111111111111" when X = 74 AND Y = 97 else
"111111111111" when X = 75 AND Y = 97 else
"111111111111" when X = 76 AND Y = 97 else
"111111111111" when X = 77 AND Y = 97 else
"111111111111" when X = 78 AND Y = 97 else
"111111111111" when X = 79 AND Y = 97 else
"111111111111" when X = 80 AND Y = 97 else
"111111111111" when X = 81 AND Y = 97 else
"111111111111" when X = 82 AND Y = 97 else
"111111111111" when X = 83 AND Y = 97 else
"111111111111" when X = 84 AND Y = 97 else
"111111111111" when X = 85 AND Y = 97 else
"111111111111" when X = 86 AND Y = 97 else
"111111111111" when X = 87 AND Y = 97 else
"111111111111" when X = 88 AND Y = 97 else
"111111111111" when X = 89 AND Y = 97 else
"111111111111" when X = 90 AND Y = 97 else
"111111111111" when X = 91 AND Y = 97 else
"111111111111" when X = 92 AND Y = 97 else
"111111111111" when X = 93 AND Y = 97 else
"111111111111" when X = 94 AND Y = 97 else
"111111111111" when X = 95 AND Y = 97 else
"111111111111" when X = 96 AND Y = 97 else
"111111111111" when X = 97 AND Y = 97 else
"111111111111" when X = 98 AND Y = 97 else
"111111111111" when X = 99 AND Y = 97 else
"111111111111" when X = 100 AND Y = 97 else
"111111111111" when X = 101 AND Y = 97 else
"111111111111" when X = 102 AND Y = 97 else
"111111111111" when X = 103 AND Y = 97 else
"111111111111" when X = 104 AND Y = 97 else
"111111111111" when X = 105 AND Y = 97 else
"111111111111" when X = 106 AND Y = 97 else
"111111111111" when X = 107 AND Y = 97 else
"111111111111" when X = 108 AND Y = 97 else
"111111111111" when X = 109 AND Y = 97 else
"111111111111" when X = 110 AND Y = 97 else
"111111111111" when X = 111 AND Y = 97 else
"111111111111" when X = 112 AND Y = 97 else
"111111111111" when X = 113 AND Y = 97 else
"111111111111" when X = 114 AND Y = 97 else
"111111111111" when X = 115 AND Y = 97 else
"111111111111" when X = 116 AND Y = 97 else
"111111111111" when X = 117 AND Y = 97 else
"111111111111" when X = 118 AND Y = 97 else
"111111111111" when X = 119 AND Y = 97 else
"111111111111" when X = 120 AND Y = 97 else
"111111111111" when X = 121 AND Y = 97 else
"111111111111" when X = 122 AND Y = 97 else
"111111111111" when X = 123 AND Y = 97 else
"111111111111" when X = 124 AND Y = 97 else
"111111111111" when X = 125 AND Y = 97 else
"111111111111" when X = 126 AND Y = 97 else
"111111111111" when X = 127 AND Y = 97 else
"111111111111" when X = 128 AND Y = 97 else
"111111111111" when X = 129 AND Y = 97 else
"111111111111" when X = 130 AND Y = 97 else
"111111111111" when X = 131 AND Y = 97 else
"111111111111" when X = 132 AND Y = 97 else
"111111111111" when X = 133 AND Y = 97 else
"111111111111" when X = 134 AND Y = 97 else
"111111111111" when X = 135 AND Y = 97 else
"111111111111" when X = 136 AND Y = 97 else
"111111111111" when X = 137 AND Y = 97 else
"111111111111" when X = 138 AND Y = 97 else
"111111111111" when X = 139 AND Y = 97 else
"111111111111" when X = 140 AND Y = 97 else
"111111111111" when X = 141 AND Y = 97 else
"111111111111" when X = 142 AND Y = 97 else
"111111111111" when X = 143 AND Y = 97 else
"111111111111" when X = 144 AND Y = 97 else
"111111111111" when X = 145 AND Y = 97 else
"111111111111" when X = 146 AND Y = 97 else
"111111111111" when X = 147 AND Y = 97 else
"111111111111" when X = 148 AND Y = 97 else
"111111111111" when X = 149 AND Y = 97 else
"111111111111" when X = 150 AND Y = 97 else
"111111111111" when X = 151 AND Y = 97 else
"111111111111" when X = 152 AND Y = 97 else
"111111111111" when X = 153 AND Y = 97 else
"111111111111" when X = 154 AND Y = 97 else
"111111111111" when X = 155 AND Y = 97 else
"111111111111" when X = 156 AND Y = 97 else
"111111111111" when X = 157 AND Y = 97 else
"111111111111" when X = 158 AND Y = 97 else
"111111111111" when X = 159 AND Y = 97 else
"111111111111" when X = 160 AND Y = 97 else
"111111111111" when X = 161 AND Y = 97 else
"111111111111" when X = 162 AND Y = 97 else
"111111111111" when X = 163 AND Y = 97 else
"111111111111" when X = 164 AND Y = 97 else
"111111111111" when X = 165 AND Y = 97 else
"111111111111" when X = 166 AND Y = 97 else
"111111111111" when X = 167 AND Y = 97 else
"111111111111" when X = 168 AND Y = 97 else
"111111111111" when X = 169 AND Y = 97 else
"111111111111" when X = 170 AND Y = 97 else
"111111111111" when X = 171 AND Y = 97 else
"111111111111" when X = 172 AND Y = 97 else
"111111111111" when X = 173 AND Y = 97 else
"111111111111" when X = 174 AND Y = 97 else
"111111111111" when X = 175 AND Y = 97 else
"111111111111" when X = 176 AND Y = 97 else
"111111111111" when X = 177 AND Y = 97 else
"111111111111" when X = 178 AND Y = 97 else
"111111111111" when X = 179 AND Y = 97 else
"111111111111" when X = 180 AND Y = 97 else
"111111111111" when X = 181 AND Y = 97 else
"111111111111" when X = 182 AND Y = 97 else
"111111111111" when X = 183 AND Y = 97 else
"111111111111" when X = 184 AND Y = 97 else
"111111111111" when X = 185 AND Y = 97 else
"111111111111" when X = 186 AND Y = 97 else
"111111111111" when X = 187 AND Y = 97 else
"111111111111" when X = 188 AND Y = 97 else
"111111111111" when X = 189 AND Y = 97 else
"111111111111" when X = 190 AND Y = 97 else
"111111111111" when X = 191 AND Y = 97 else
"111111111111" when X = 192 AND Y = 97 else
"111111111111" when X = 193 AND Y = 97 else
"111111111111" when X = 194 AND Y = 97 else
"111111111111" when X = 195 AND Y = 97 else
"111111111111" when X = 196 AND Y = 97 else
"111111111111" when X = 197 AND Y = 97 else
"111111111111" when X = 198 AND Y = 97 else
"111111111111" when X = 199 AND Y = 97 else
"111111111111" when X = 200 AND Y = 97 else
"111111111111" when X = 201 AND Y = 97 else
"111111111111" when X = 202 AND Y = 97 else
"111111111111" when X = 203 AND Y = 97 else
"111111111111" when X = 204 AND Y = 97 else
"110111011111" when X = 205 AND Y = 97 else
"110111011111" when X = 206 AND Y = 97 else
"110111011111" when X = 207 AND Y = 97 else
"110111011111" when X = 208 AND Y = 97 else
"110111011111" when X = 209 AND Y = 97 else
"110111011111" when X = 210 AND Y = 97 else
"110111011111" when X = 211 AND Y = 97 else
"110111011111" when X = 212 AND Y = 97 else
"110111011111" when X = 213 AND Y = 97 else
"110111011111" when X = 214 AND Y = 97 else
"110111011111" when X = 215 AND Y = 97 else
"110111011111" when X = 216 AND Y = 97 else
"110111011111" when X = 217 AND Y = 97 else
"110111011111" when X = 218 AND Y = 97 else
"110111011111" when X = 219 AND Y = 97 else
"111111111111" when X = 220 AND Y = 97 else
"111111111111" when X = 221 AND Y = 97 else
"111111111111" when X = 222 AND Y = 97 else
"111111111111" when X = 223 AND Y = 97 else
"111111111111" when X = 224 AND Y = 97 else
"111111111111" when X = 225 AND Y = 97 else
"111111111111" when X = 226 AND Y = 97 else
"111111111111" when X = 227 AND Y = 97 else
"111111111111" when X = 228 AND Y = 97 else
"111111111111" when X = 229 AND Y = 97 else
"111111111111" when X = 230 AND Y = 97 else
"111111111111" when X = 231 AND Y = 97 else
"111111111111" when X = 232 AND Y = 97 else
"111111111111" when X = 233 AND Y = 97 else
"111111111111" when X = 234 AND Y = 97 else
"111111111111" when X = 235 AND Y = 97 else
"111111111111" when X = 236 AND Y = 97 else
"111111111111" when X = 237 AND Y = 97 else
"111111111111" when X = 238 AND Y = 97 else
"111111111111" when X = 239 AND Y = 97 else
"111111111111" when X = 240 AND Y = 97 else
"111111111111" when X = 241 AND Y = 97 else
"111111111111" when X = 242 AND Y = 97 else
"111111111111" when X = 243 AND Y = 97 else
"111111111111" when X = 244 AND Y = 97 else
"111111111111" when X = 245 AND Y = 97 else
"111111111111" when X = 246 AND Y = 97 else
"111111111111" when X = 247 AND Y = 97 else
"111111111111" when X = 248 AND Y = 97 else
"111111111111" when X = 249 AND Y = 97 else
"111111111111" when X = 250 AND Y = 97 else
"111111111111" when X = 251 AND Y = 97 else
"111111111111" when X = 252 AND Y = 97 else
"111111111111" when X = 253 AND Y = 97 else
"111111111111" when X = 254 AND Y = 97 else
"111111111111" when X = 255 AND Y = 97 else
"111111111111" when X = 256 AND Y = 97 else
"111111111111" when X = 257 AND Y = 97 else
"111111111111" when X = 258 AND Y = 97 else
"111111111111" when X = 259 AND Y = 97 else
"111111111111" when X = 260 AND Y = 97 else
"111111111111" when X = 261 AND Y = 97 else
"111111111111" when X = 262 AND Y = 97 else
"111111111111" when X = 263 AND Y = 97 else
"111111111111" when X = 264 AND Y = 97 else
"111111111111" when X = 265 AND Y = 97 else
"111111111111" when X = 266 AND Y = 97 else
"111111111111" when X = 267 AND Y = 97 else
"111111111111" when X = 268 AND Y = 97 else
"111111111111" when X = 269 AND Y = 97 else
"111111111111" when X = 270 AND Y = 97 else
"111111111111" when X = 271 AND Y = 97 else
"111111111111" when X = 272 AND Y = 97 else
"111111111111" when X = 273 AND Y = 97 else
"111111111111" when X = 274 AND Y = 97 else
"110111011111" when X = 275 AND Y = 97 else
"110111011111" when X = 276 AND Y = 97 else
"110111011111" when X = 277 AND Y = 97 else
"110111011111" when X = 278 AND Y = 97 else
"110111011111" when X = 279 AND Y = 97 else
"110111011111" when X = 280 AND Y = 97 else
"110111011111" when X = 281 AND Y = 97 else
"110111011111" when X = 282 AND Y = 97 else
"110111011111" when X = 283 AND Y = 97 else
"110111011111" when X = 284 AND Y = 97 else
"111111111111" when X = 285 AND Y = 97 else
"111111111111" when X = 286 AND Y = 97 else
"111111111111" when X = 287 AND Y = 97 else
"111111111111" when X = 288 AND Y = 97 else
"111111111111" when X = 289 AND Y = 97 else
"111111111111" when X = 290 AND Y = 97 else
"111111111111" when X = 291 AND Y = 97 else
"111111111111" when X = 292 AND Y = 97 else
"111111111111" when X = 293 AND Y = 97 else
"111111111111" when X = 294 AND Y = 97 else
"111111111111" when X = 295 AND Y = 97 else
"111111111111" when X = 296 AND Y = 97 else
"111111111111" when X = 297 AND Y = 97 else
"111111111111" when X = 298 AND Y = 97 else
"111111111111" when X = 299 AND Y = 97 else
"111111111111" when X = 300 AND Y = 97 else
"111111111111" when X = 301 AND Y = 97 else
"111111111111" when X = 302 AND Y = 97 else
"111111111111" when X = 303 AND Y = 97 else
"111111111111" when X = 304 AND Y = 97 else
"110111011111" when X = 305 AND Y = 97 else
"110111011111" when X = 306 AND Y = 97 else
"110111011111" when X = 307 AND Y = 97 else
"110111011111" when X = 308 AND Y = 97 else
"110111011111" when X = 309 AND Y = 97 else
"110111011111" when X = 310 AND Y = 97 else
"110111011111" when X = 311 AND Y = 97 else
"110111011111" when X = 312 AND Y = 97 else
"110111011111" when X = 313 AND Y = 97 else
"110111011111" when X = 314 AND Y = 97 else
"110111011111" when X = 315 AND Y = 97 else
"110111011111" when X = 316 AND Y = 97 else
"110111011111" when X = 317 AND Y = 97 else
"110111011111" when X = 318 AND Y = 97 else
"110111011111" when X = 319 AND Y = 97 else
"110111011111" when X = 320 AND Y = 97 else
"110111011111" when X = 321 AND Y = 97 else
"110111011111" when X = 322 AND Y = 97 else
"110111011111" when X = 323 AND Y = 97 else
"110111011111" when X = 324 AND Y = 97 else
"100010011101" when X = 0 AND Y = 98 else
"100010011101" when X = 1 AND Y = 98 else
"100010011101" when X = 2 AND Y = 98 else
"100010011101" when X = 3 AND Y = 98 else
"100010011101" when X = 4 AND Y = 98 else
"100010011101" when X = 5 AND Y = 98 else
"100010011101" when X = 6 AND Y = 98 else
"100010011101" when X = 7 AND Y = 98 else
"100010011101" when X = 8 AND Y = 98 else
"100010011101" when X = 9 AND Y = 98 else
"100010011101" when X = 10 AND Y = 98 else
"100010011101" when X = 11 AND Y = 98 else
"100010011101" when X = 12 AND Y = 98 else
"100010011101" when X = 13 AND Y = 98 else
"100010011101" when X = 14 AND Y = 98 else
"110111011111" when X = 15 AND Y = 98 else
"110111011111" when X = 16 AND Y = 98 else
"110111011111" when X = 17 AND Y = 98 else
"110111011111" when X = 18 AND Y = 98 else
"110111011111" when X = 19 AND Y = 98 else
"110111011111" when X = 20 AND Y = 98 else
"110111011111" when X = 21 AND Y = 98 else
"110111011111" when X = 22 AND Y = 98 else
"110111011111" when X = 23 AND Y = 98 else
"110111011111" when X = 24 AND Y = 98 else
"110111011111" when X = 25 AND Y = 98 else
"110111011111" when X = 26 AND Y = 98 else
"110111011111" when X = 27 AND Y = 98 else
"110111011111" when X = 28 AND Y = 98 else
"110111011111" when X = 29 AND Y = 98 else
"110111011111" when X = 30 AND Y = 98 else
"110111011111" when X = 31 AND Y = 98 else
"110111011111" when X = 32 AND Y = 98 else
"110111011111" when X = 33 AND Y = 98 else
"110111011111" when X = 34 AND Y = 98 else
"110111011111" when X = 35 AND Y = 98 else
"110111011111" when X = 36 AND Y = 98 else
"110111011111" when X = 37 AND Y = 98 else
"110111011111" when X = 38 AND Y = 98 else
"110111011111" when X = 39 AND Y = 98 else
"110111011111" when X = 40 AND Y = 98 else
"110111011111" when X = 41 AND Y = 98 else
"110111011111" when X = 42 AND Y = 98 else
"110111011111" when X = 43 AND Y = 98 else
"110111011111" when X = 44 AND Y = 98 else
"110111011111" when X = 45 AND Y = 98 else
"110111011111" when X = 46 AND Y = 98 else
"110111011111" when X = 47 AND Y = 98 else
"110111011111" when X = 48 AND Y = 98 else
"110111011111" when X = 49 AND Y = 98 else
"110111011111" when X = 50 AND Y = 98 else
"110111011111" when X = 51 AND Y = 98 else
"110111011111" when X = 52 AND Y = 98 else
"110111011111" when X = 53 AND Y = 98 else
"110111011111" when X = 54 AND Y = 98 else
"110111011111" when X = 55 AND Y = 98 else
"110111011111" when X = 56 AND Y = 98 else
"110111011111" when X = 57 AND Y = 98 else
"110111011111" when X = 58 AND Y = 98 else
"110111011111" when X = 59 AND Y = 98 else
"110111011111" when X = 60 AND Y = 98 else
"110111011111" when X = 61 AND Y = 98 else
"110111011111" when X = 62 AND Y = 98 else
"110111011111" when X = 63 AND Y = 98 else
"110111011111" when X = 64 AND Y = 98 else
"110111011111" when X = 65 AND Y = 98 else
"110111011111" when X = 66 AND Y = 98 else
"110111011111" when X = 67 AND Y = 98 else
"110111011111" when X = 68 AND Y = 98 else
"110111011111" when X = 69 AND Y = 98 else
"111111111111" when X = 70 AND Y = 98 else
"111111111111" when X = 71 AND Y = 98 else
"111111111111" when X = 72 AND Y = 98 else
"111111111111" when X = 73 AND Y = 98 else
"111111111111" when X = 74 AND Y = 98 else
"111111111111" when X = 75 AND Y = 98 else
"111111111111" when X = 76 AND Y = 98 else
"111111111111" when X = 77 AND Y = 98 else
"111111111111" when X = 78 AND Y = 98 else
"111111111111" when X = 79 AND Y = 98 else
"111111111111" when X = 80 AND Y = 98 else
"111111111111" when X = 81 AND Y = 98 else
"111111111111" when X = 82 AND Y = 98 else
"111111111111" when X = 83 AND Y = 98 else
"111111111111" when X = 84 AND Y = 98 else
"111111111111" when X = 85 AND Y = 98 else
"111111111111" when X = 86 AND Y = 98 else
"111111111111" when X = 87 AND Y = 98 else
"111111111111" when X = 88 AND Y = 98 else
"111111111111" when X = 89 AND Y = 98 else
"111111111111" when X = 90 AND Y = 98 else
"111111111111" when X = 91 AND Y = 98 else
"111111111111" when X = 92 AND Y = 98 else
"111111111111" when X = 93 AND Y = 98 else
"111111111111" when X = 94 AND Y = 98 else
"111111111111" when X = 95 AND Y = 98 else
"111111111111" when X = 96 AND Y = 98 else
"111111111111" when X = 97 AND Y = 98 else
"111111111111" when X = 98 AND Y = 98 else
"111111111111" when X = 99 AND Y = 98 else
"111111111111" when X = 100 AND Y = 98 else
"111111111111" when X = 101 AND Y = 98 else
"111111111111" when X = 102 AND Y = 98 else
"111111111111" when X = 103 AND Y = 98 else
"111111111111" when X = 104 AND Y = 98 else
"111111111111" when X = 105 AND Y = 98 else
"111111111111" when X = 106 AND Y = 98 else
"111111111111" when X = 107 AND Y = 98 else
"111111111111" when X = 108 AND Y = 98 else
"111111111111" when X = 109 AND Y = 98 else
"111111111111" when X = 110 AND Y = 98 else
"111111111111" when X = 111 AND Y = 98 else
"111111111111" when X = 112 AND Y = 98 else
"111111111111" when X = 113 AND Y = 98 else
"111111111111" when X = 114 AND Y = 98 else
"111111111111" when X = 115 AND Y = 98 else
"111111111111" when X = 116 AND Y = 98 else
"111111111111" when X = 117 AND Y = 98 else
"111111111111" when X = 118 AND Y = 98 else
"111111111111" when X = 119 AND Y = 98 else
"111111111111" when X = 120 AND Y = 98 else
"111111111111" when X = 121 AND Y = 98 else
"111111111111" when X = 122 AND Y = 98 else
"111111111111" when X = 123 AND Y = 98 else
"111111111111" when X = 124 AND Y = 98 else
"111111111111" when X = 125 AND Y = 98 else
"111111111111" when X = 126 AND Y = 98 else
"111111111111" when X = 127 AND Y = 98 else
"111111111111" when X = 128 AND Y = 98 else
"111111111111" when X = 129 AND Y = 98 else
"111111111111" when X = 130 AND Y = 98 else
"111111111111" when X = 131 AND Y = 98 else
"111111111111" when X = 132 AND Y = 98 else
"111111111111" when X = 133 AND Y = 98 else
"111111111111" when X = 134 AND Y = 98 else
"111111111111" when X = 135 AND Y = 98 else
"111111111111" when X = 136 AND Y = 98 else
"111111111111" when X = 137 AND Y = 98 else
"111111111111" when X = 138 AND Y = 98 else
"111111111111" when X = 139 AND Y = 98 else
"111111111111" when X = 140 AND Y = 98 else
"111111111111" when X = 141 AND Y = 98 else
"111111111111" when X = 142 AND Y = 98 else
"111111111111" when X = 143 AND Y = 98 else
"111111111111" when X = 144 AND Y = 98 else
"111111111111" when X = 145 AND Y = 98 else
"111111111111" when X = 146 AND Y = 98 else
"111111111111" when X = 147 AND Y = 98 else
"111111111111" when X = 148 AND Y = 98 else
"111111111111" when X = 149 AND Y = 98 else
"111111111111" when X = 150 AND Y = 98 else
"111111111111" when X = 151 AND Y = 98 else
"111111111111" when X = 152 AND Y = 98 else
"111111111111" when X = 153 AND Y = 98 else
"111111111111" when X = 154 AND Y = 98 else
"111111111111" when X = 155 AND Y = 98 else
"111111111111" when X = 156 AND Y = 98 else
"111111111111" when X = 157 AND Y = 98 else
"111111111111" when X = 158 AND Y = 98 else
"111111111111" when X = 159 AND Y = 98 else
"111111111111" when X = 160 AND Y = 98 else
"111111111111" when X = 161 AND Y = 98 else
"111111111111" when X = 162 AND Y = 98 else
"111111111111" when X = 163 AND Y = 98 else
"111111111111" when X = 164 AND Y = 98 else
"111111111111" when X = 165 AND Y = 98 else
"111111111111" when X = 166 AND Y = 98 else
"111111111111" when X = 167 AND Y = 98 else
"111111111111" when X = 168 AND Y = 98 else
"111111111111" when X = 169 AND Y = 98 else
"111111111111" when X = 170 AND Y = 98 else
"111111111111" when X = 171 AND Y = 98 else
"111111111111" when X = 172 AND Y = 98 else
"111111111111" when X = 173 AND Y = 98 else
"111111111111" when X = 174 AND Y = 98 else
"111111111111" when X = 175 AND Y = 98 else
"111111111111" when X = 176 AND Y = 98 else
"111111111111" when X = 177 AND Y = 98 else
"111111111111" when X = 178 AND Y = 98 else
"111111111111" when X = 179 AND Y = 98 else
"111111111111" when X = 180 AND Y = 98 else
"111111111111" when X = 181 AND Y = 98 else
"111111111111" when X = 182 AND Y = 98 else
"111111111111" when X = 183 AND Y = 98 else
"111111111111" when X = 184 AND Y = 98 else
"111111111111" when X = 185 AND Y = 98 else
"111111111111" when X = 186 AND Y = 98 else
"111111111111" when X = 187 AND Y = 98 else
"111111111111" when X = 188 AND Y = 98 else
"111111111111" when X = 189 AND Y = 98 else
"111111111111" when X = 190 AND Y = 98 else
"111111111111" when X = 191 AND Y = 98 else
"111111111111" when X = 192 AND Y = 98 else
"111111111111" when X = 193 AND Y = 98 else
"111111111111" when X = 194 AND Y = 98 else
"111111111111" when X = 195 AND Y = 98 else
"111111111111" when X = 196 AND Y = 98 else
"111111111111" when X = 197 AND Y = 98 else
"111111111111" when X = 198 AND Y = 98 else
"111111111111" when X = 199 AND Y = 98 else
"111111111111" when X = 200 AND Y = 98 else
"111111111111" when X = 201 AND Y = 98 else
"111111111111" when X = 202 AND Y = 98 else
"111111111111" when X = 203 AND Y = 98 else
"111111111111" when X = 204 AND Y = 98 else
"110111011111" when X = 205 AND Y = 98 else
"110111011111" when X = 206 AND Y = 98 else
"110111011111" when X = 207 AND Y = 98 else
"110111011111" when X = 208 AND Y = 98 else
"110111011111" when X = 209 AND Y = 98 else
"110111011111" when X = 210 AND Y = 98 else
"110111011111" when X = 211 AND Y = 98 else
"110111011111" when X = 212 AND Y = 98 else
"110111011111" when X = 213 AND Y = 98 else
"110111011111" when X = 214 AND Y = 98 else
"110111011111" when X = 215 AND Y = 98 else
"110111011111" when X = 216 AND Y = 98 else
"110111011111" when X = 217 AND Y = 98 else
"110111011111" when X = 218 AND Y = 98 else
"110111011111" when X = 219 AND Y = 98 else
"111111111111" when X = 220 AND Y = 98 else
"111111111111" when X = 221 AND Y = 98 else
"111111111111" when X = 222 AND Y = 98 else
"111111111111" when X = 223 AND Y = 98 else
"111111111111" when X = 224 AND Y = 98 else
"111111111111" when X = 225 AND Y = 98 else
"111111111111" when X = 226 AND Y = 98 else
"111111111111" when X = 227 AND Y = 98 else
"111111111111" when X = 228 AND Y = 98 else
"111111111111" when X = 229 AND Y = 98 else
"111111111111" when X = 230 AND Y = 98 else
"111111111111" when X = 231 AND Y = 98 else
"111111111111" when X = 232 AND Y = 98 else
"111111111111" when X = 233 AND Y = 98 else
"111111111111" when X = 234 AND Y = 98 else
"111111111111" when X = 235 AND Y = 98 else
"111111111111" when X = 236 AND Y = 98 else
"111111111111" when X = 237 AND Y = 98 else
"111111111111" when X = 238 AND Y = 98 else
"111111111111" when X = 239 AND Y = 98 else
"111111111111" when X = 240 AND Y = 98 else
"111111111111" when X = 241 AND Y = 98 else
"111111111111" when X = 242 AND Y = 98 else
"111111111111" when X = 243 AND Y = 98 else
"111111111111" when X = 244 AND Y = 98 else
"111111111111" when X = 245 AND Y = 98 else
"111111111111" when X = 246 AND Y = 98 else
"111111111111" when X = 247 AND Y = 98 else
"111111111111" when X = 248 AND Y = 98 else
"111111111111" when X = 249 AND Y = 98 else
"111111111111" when X = 250 AND Y = 98 else
"111111111111" when X = 251 AND Y = 98 else
"111111111111" when X = 252 AND Y = 98 else
"111111111111" when X = 253 AND Y = 98 else
"111111111111" when X = 254 AND Y = 98 else
"111111111111" when X = 255 AND Y = 98 else
"111111111111" when X = 256 AND Y = 98 else
"111111111111" when X = 257 AND Y = 98 else
"111111111111" when X = 258 AND Y = 98 else
"111111111111" when X = 259 AND Y = 98 else
"111111111111" when X = 260 AND Y = 98 else
"111111111111" when X = 261 AND Y = 98 else
"111111111111" when X = 262 AND Y = 98 else
"111111111111" when X = 263 AND Y = 98 else
"111111111111" when X = 264 AND Y = 98 else
"111111111111" when X = 265 AND Y = 98 else
"111111111111" when X = 266 AND Y = 98 else
"111111111111" when X = 267 AND Y = 98 else
"111111111111" when X = 268 AND Y = 98 else
"111111111111" when X = 269 AND Y = 98 else
"111111111111" when X = 270 AND Y = 98 else
"111111111111" when X = 271 AND Y = 98 else
"111111111111" when X = 272 AND Y = 98 else
"111111111111" when X = 273 AND Y = 98 else
"111111111111" when X = 274 AND Y = 98 else
"110111011111" when X = 275 AND Y = 98 else
"110111011111" when X = 276 AND Y = 98 else
"110111011111" when X = 277 AND Y = 98 else
"110111011111" when X = 278 AND Y = 98 else
"110111011111" when X = 279 AND Y = 98 else
"110111011111" when X = 280 AND Y = 98 else
"110111011111" when X = 281 AND Y = 98 else
"110111011111" when X = 282 AND Y = 98 else
"110111011111" when X = 283 AND Y = 98 else
"110111011111" when X = 284 AND Y = 98 else
"111111111111" when X = 285 AND Y = 98 else
"111111111111" when X = 286 AND Y = 98 else
"111111111111" when X = 287 AND Y = 98 else
"111111111111" when X = 288 AND Y = 98 else
"111111111111" when X = 289 AND Y = 98 else
"111111111111" when X = 290 AND Y = 98 else
"111111111111" when X = 291 AND Y = 98 else
"111111111111" when X = 292 AND Y = 98 else
"111111111111" when X = 293 AND Y = 98 else
"111111111111" when X = 294 AND Y = 98 else
"111111111111" when X = 295 AND Y = 98 else
"111111111111" when X = 296 AND Y = 98 else
"111111111111" when X = 297 AND Y = 98 else
"111111111111" when X = 298 AND Y = 98 else
"111111111111" when X = 299 AND Y = 98 else
"111111111111" when X = 300 AND Y = 98 else
"111111111111" when X = 301 AND Y = 98 else
"111111111111" when X = 302 AND Y = 98 else
"111111111111" when X = 303 AND Y = 98 else
"111111111111" when X = 304 AND Y = 98 else
"110111011111" when X = 305 AND Y = 98 else
"110111011111" when X = 306 AND Y = 98 else
"110111011111" when X = 307 AND Y = 98 else
"110111011111" when X = 308 AND Y = 98 else
"110111011111" when X = 309 AND Y = 98 else
"110111011111" when X = 310 AND Y = 98 else
"110111011111" when X = 311 AND Y = 98 else
"110111011111" when X = 312 AND Y = 98 else
"110111011111" when X = 313 AND Y = 98 else
"110111011111" when X = 314 AND Y = 98 else
"110111011111" when X = 315 AND Y = 98 else
"110111011111" when X = 316 AND Y = 98 else
"110111011111" when X = 317 AND Y = 98 else
"110111011111" when X = 318 AND Y = 98 else
"110111011111" when X = 319 AND Y = 98 else
"110111011111" when X = 320 AND Y = 98 else
"110111011111" when X = 321 AND Y = 98 else
"110111011111" when X = 322 AND Y = 98 else
"110111011111" when X = 323 AND Y = 98 else
"110111011111" when X = 324 AND Y = 98 else
"100010011101" when X = 0 AND Y = 99 else
"100010011101" when X = 1 AND Y = 99 else
"100010011101" when X = 2 AND Y = 99 else
"100010011101" when X = 3 AND Y = 99 else
"100010011101" when X = 4 AND Y = 99 else
"100010011101" when X = 5 AND Y = 99 else
"100010011101" when X = 6 AND Y = 99 else
"100010011101" when X = 7 AND Y = 99 else
"100010011101" when X = 8 AND Y = 99 else
"100010011101" when X = 9 AND Y = 99 else
"100010011101" when X = 10 AND Y = 99 else
"100010011101" when X = 11 AND Y = 99 else
"100010011101" when X = 12 AND Y = 99 else
"100010011101" when X = 13 AND Y = 99 else
"100010011101" when X = 14 AND Y = 99 else
"110111011111" when X = 15 AND Y = 99 else
"110111011111" when X = 16 AND Y = 99 else
"110111011111" when X = 17 AND Y = 99 else
"110111011111" when X = 18 AND Y = 99 else
"110111011111" when X = 19 AND Y = 99 else
"110111011111" when X = 20 AND Y = 99 else
"110111011111" when X = 21 AND Y = 99 else
"110111011111" when X = 22 AND Y = 99 else
"110111011111" when X = 23 AND Y = 99 else
"110111011111" when X = 24 AND Y = 99 else
"110111011111" when X = 25 AND Y = 99 else
"110111011111" when X = 26 AND Y = 99 else
"110111011111" when X = 27 AND Y = 99 else
"110111011111" when X = 28 AND Y = 99 else
"110111011111" when X = 29 AND Y = 99 else
"110111011111" when X = 30 AND Y = 99 else
"110111011111" when X = 31 AND Y = 99 else
"110111011111" when X = 32 AND Y = 99 else
"110111011111" when X = 33 AND Y = 99 else
"110111011111" when X = 34 AND Y = 99 else
"110111011111" when X = 35 AND Y = 99 else
"110111011111" when X = 36 AND Y = 99 else
"110111011111" when X = 37 AND Y = 99 else
"110111011111" when X = 38 AND Y = 99 else
"110111011111" when X = 39 AND Y = 99 else
"110111011111" when X = 40 AND Y = 99 else
"110111011111" when X = 41 AND Y = 99 else
"110111011111" when X = 42 AND Y = 99 else
"110111011111" when X = 43 AND Y = 99 else
"110111011111" when X = 44 AND Y = 99 else
"110111011111" when X = 45 AND Y = 99 else
"110111011111" when X = 46 AND Y = 99 else
"110111011111" when X = 47 AND Y = 99 else
"110111011111" when X = 48 AND Y = 99 else
"110111011111" when X = 49 AND Y = 99 else
"110111011111" when X = 50 AND Y = 99 else
"110111011111" when X = 51 AND Y = 99 else
"110111011111" when X = 52 AND Y = 99 else
"110111011111" when X = 53 AND Y = 99 else
"110111011111" when X = 54 AND Y = 99 else
"110111011111" when X = 55 AND Y = 99 else
"110111011111" when X = 56 AND Y = 99 else
"110111011111" when X = 57 AND Y = 99 else
"110111011111" when X = 58 AND Y = 99 else
"110111011111" when X = 59 AND Y = 99 else
"110111011111" when X = 60 AND Y = 99 else
"110111011111" when X = 61 AND Y = 99 else
"110111011111" when X = 62 AND Y = 99 else
"110111011111" when X = 63 AND Y = 99 else
"110111011111" when X = 64 AND Y = 99 else
"110111011111" when X = 65 AND Y = 99 else
"110111011111" when X = 66 AND Y = 99 else
"110111011111" when X = 67 AND Y = 99 else
"110111011111" when X = 68 AND Y = 99 else
"110111011111" when X = 69 AND Y = 99 else
"111111111111" when X = 70 AND Y = 99 else
"111111111111" when X = 71 AND Y = 99 else
"111111111111" when X = 72 AND Y = 99 else
"111111111111" when X = 73 AND Y = 99 else
"111111111111" when X = 74 AND Y = 99 else
"111111111111" when X = 75 AND Y = 99 else
"111111111111" when X = 76 AND Y = 99 else
"111111111111" when X = 77 AND Y = 99 else
"111111111111" when X = 78 AND Y = 99 else
"111111111111" when X = 79 AND Y = 99 else
"111111111111" when X = 80 AND Y = 99 else
"111111111111" when X = 81 AND Y = 99 else
"111111111111" when X = 82 AND Y = 99 else
"111111111111" when X = 83 AND Y = 99 else
"111111111111" when X = 84 AND Y = 99 else
"111111111111" when X = 85 AND Y = 99 else
"111111111111" when X = 86 AND Y = 99 else
"111111111111" when X = 87 AND Y = 99 else
"111111111111" when X = 88 AND Y = 99 else
"111111111111" when X = 89 AND Y = 99 else
"111111111111" when X = 90 AND Y = 99 else
"111111111111" when X = 91 AND Y = 99 else
"111111111111" when X = 92 AND Y = 99 else
"111111111111" when X = 93 AND Y = 99 else
"111111111111" when X = 94 AND Y = 99 else
"111111111111" when X = 95 AND Y = 99 else
"111111111111" when X = 96 AND Y = 99 else
"111111111111" when X = 97 AND Y = 99 else
"111111111111" when X = 98 AND Y = 99 else
"111111111111" when X = 99 AND Y = 99 else
"111111111111" when X = 100 AND Y = 99 else
"111111111111" when X = 101 AND Y = 99 else
"111111111111" when X = 102 AND Y = 99 else
"111111111111" when X = 103 AND Y = 99 else
"111111111111" when X = 104 AND Y = 99 else
"111111111111" when X = 105 AND Y = 99 else
"111111111111" when X = 106 AND Y = 99 else
"111111111111" when X = 107 AND Y = 99 else
"111111111111" when X = 108 AND Y = 99 else
"111111111111" when X = 109 AND Y = 99 else
"111111111111" when X = 110 AND Y = 99 else
"111111111111" when X = 111 AND Y = 99 else
"111111111111" when X = 112 AND Y = 99 else
"111111111111" when X = 113 AND Y = 99 else
"111111111111" when X = 114 AND Y = 99 else
"111111111111" when X = 115 AND Y = 99 else
"111111111111" when X = 116 AND Y = 99 else
"111111111111" when X = 117 AND Y = 99 else
"111111111111" when X = 118 AND Y = 99 else
"111111111111" when X = 119 AND Y = 99 else
"111111111111" when X = 120 AND Y = 99 else
"111111111111" when X = 121 AND Y = 99 else
"111111111111" when X = 122 AND Y = 99 else
"111111111111" when X = 123 AND Y = 99 else
"111111111111" when X = 124 AND Y = 99 else
"111111111111" when X = 125 AND Y = 99 else
"111111111111" when X = 126 AND Y = 99 else
"111111111111" when X = 127 AND Y = 99 else
"111111111111" when X = 128 AND Y = 99 else
"111111111111" when X = 129 AND Y = 99 else
"111111111111" when X = 130 AND Y = 99 else
"111111111111" when X = 131 AND Y = 99 else
"111111111111" when X = 132 AND Y = 99 else
"111111111111" when X = 133 AND Y = 99 else
"111111111111" when X = 134 AND Y = 99 else
"111111111111" when X = 135 AND Y = 99 else
"111111111111" when X = 136 AND Y = 99 else
"111111111111" when X = 137 AND Y = 99 else
"111111111111" when X = 138 AND Y = 99 else
"111111111111" when X = 139 AND Y = 99 else
"111111111111" when X = 140 AND Y = 99 else
"111111111111" when X = 141 AND Y = 99 else
"111111111111" when X = 142 AND Y = 99 else
"111111111111" when X = 143 AND Y = 99 else
"111111111111" when X = 144 AND Y = 99 else
"111111111111" when X = 145 AND Y = 99 else
"111111111111" when X = 146 AND Y = 99 else
"111111111111" when X = 147 AND Y = 99 else
"111111111111" when X = 148 AND Y = 99 else
"111111111111" when X = 149 AND Y = 99 else
"111111111111" when X = 150 AND Y = 99 else
"111111111111" when X = 151 AND Y = 99 else
"111111111111" when X = 152 AND Y = 99 else
"111111111111" when X = 153 AND Y = 99 else
"111111111111" when X = 154 AND Y = 99 else
"111111111111" when X = 155 AND Y = 99 else
"111111111111" when X = 156 AND Y = 99 else
"111111111111" when X = 157 AND Y = 99 else
"111111111111" when X = 158 AND Y = 99 else
"111111111111" when X = 159 AND Y = 99 else
"111111111111" when X = 160 AND Y = 99 else
"111111111111" when X = 161 AND Y = 99 else
"111111111111" when X = 162 AND Y = 99 else
"111111111111" when X = 163 AND Y = 99 else
"111111111111" when X = 164 AND Y = 99 else
"111111111111" when X = 165 AND Y = 99 else
"111111111111" when X = 166 AND Y = 99 else
"111111111111" when X = 167 AND Y = 99 else
"111111111111" when X = 168 AND Y = 99 else
"111111111111" when X = 169 AND Y = 99 else
"111111111111" when X = 170 AND Y = 99 else
"111111111111" when X = 171 AND Y = 99 else
"111111111111" when X = 172 AND Y = 99 else
"111111111111" when X = 173 AND Y = 99 else
"111111111111" when X = 174 AND Y = 99 else
"111111111111" when X = 175 AND Y = 99 else
"111111111111" when X = 176 AND Y = 99 else
"111111111111" when X = 177 AND Y = 99 else
"111111111111" when X = 178 AND Y = 99 else
"111111111111" when X = 179 AND Y = 99 else
"111111111111" when X = 180 AND Y = 99 else
"111111111111" when X = 181 AND Y = 99 else
"111111111111" when X = 182 AND Y = 99 else
"111111111111" when X = 183 AND Y = 99 else
"111111111111" when X = 184 AND Y = 99 else
"111111111111" when X = 185 AND Y = 99 else
"111111111111" when X = 186 AND Y = 99 else
"111111111111" when X = 187 AND Y = 99 else
"111111111111" when X = 188 AND Y = 99 else
"111111111111" when X = 189 AND Y = 99 else
"111111111111" when X = 190 AND Y = 99 else
"111111111111" when X = 191 AND Y = 99 else
"111111111111" when X = 192 AND Y = 99 else
"111111111111" when X = 193 AND Y = 99 else
"111111111111" when X = 194 AND Y = 99 else
"111111111111" when X = 195 AND Y = 99 else
"111111111111" when X = 196 AND Y = 99 else
"111111111111" when X = 197 AND Y = 99 else
"111111111111" when X = 198 AND Y = 99 else
"111111111111" when X = 199 AND Y = 99 else
"111111111111" when X = 200 AND Y = 99 else
"111111111111" when X = 201 AND Y = 99 else
"111111111111" when X = 202 AND Y = 99 else
"111111111111" when X = 203 AND Y = 99 else
"111111111111" when X = 204 AND Y = 99 else
"110111011111" when X = 205 AND Y = 99 else
"110111011111" when X = 206 AND Y = 99 else
"110111011111" when X = 207 AND Y = 99 else
"110111011111" when X = 208 AND Y = 99 else
"110111011111" when X = 209 AND Y = 99 else
"110111011111" when X = 210 AND Y = 99 else
"110111011111" when X = 211 AND Y = 99 else
"110111011111" when X = 212 AND Y = 99 else
"110111011111" when X = 213 AND Y = 99 else
"110111011111" when X = 214 AND Y = 99 else
"110111011111" when X = 215 AND Y = 99 else
"110111011111" when X = 216 AND Y = 99 else
"110111011111" when X = 217 AND Y = 99 else
"110111011111" when X = 218 AND Y = 99 else
"110111011111" when X = 219 AND Y = 99 else
"111111111111" when X = 220 AND Y = 99 else
"111111111111" when X = 221 AND Y = 99 else
"111111111111" when X = 222 AND Y = 99 else
"111111111111" when X = 223 AND Y = 99 else
"111111111111" when X = 224 AND Y = 99 else
"111111111111" when X = 225 AND Y = 99 else
"111111111111" when X = 226 AND Y = 99 else
"111111111111" when X = 227 AND Y = 99 else
"111111111111" when X = 228 AND Y = 99 else
"111111111111" when X = 229 AND Y = 99 else
"111111111111" when X = 230 AND Y = 99 else
"111111111111" when X = 231 AND Y = 99 else
"111111111111" when X = 232 AND Y = 99 else
"111111111111" when X = 233 AND Y = 99 else
"111111111111" when X = 234 AND Y = 99 else
"111111111111" when X = 235 AND Y = 99 else
"111111111111" when X = 236 AND Y = 99 else
"111111111111" when X = 237 AND Y = 99 else
"111111111111" when X = 238 AND Y = 99 else
"111111111111" when X = 239 AND Y = 99 else
"111111111111" when X = 240 AND Y = 99 else
"111111111111" when X = 241 AND Y = 99 else
"111111111111" when X = 242 AND Y = 99 else
"111111111111" when X = 243 AND Y = 99 else
"111111111111" when X = 244 AND Y = 99 else
"111111111111" when X = 245 AND Y = 99 else
"111111111111" when X = 246 AND Y = 99 else
"111111111111" when X = 247 AND Y = 99 else
"111111111111" when X = 248 AND Y = 99 else
"111111111111" when X = 249 AND Y = 99 else
"111111111111" when X = 250 AND Y = 99 else
"111111111111" when X = 251 AND Y = 99 else
"111111111111" when X = 252 AND Y = 99 else
"111111111111" when X = 253 AND Y = 99 else
"111111111111" when X = 254 AND Y = 99 else
"111111111111" when X = 255 AND Y = 99 else
"111111111111" when X = 256 AND Y = 99 else
"111111111111" when X = 257 AND Y = 99 else
"111111111111" when X = 258 AND Y = 99 else
"111111111111" when X = 259 AND Y = 99 else
"111111111111" when X = 260 AND Y = 99 else
"111111111111" when X = 261 AND Y = 99 else
"111111111111" when X = 262 AND Y = 99 else
"111111111111" when X = 263 AND Y = 99 else
"111111111111" when X = 264 AND Y = 99 else
"111111111111" when X = 265 AND Y = 99 else
"111111111111" when X = 266 AND Y = 99 else
"111111111111" when X = 267 AND Y = 99 else
"111111111111" when X = 268 AND Y = 99 else
"111111111111" when X = 269 AND Y = 99 else
"111111111111" when X = 270 AND Y = 99 else
"111111111111" when X = 271 AND Y = 99 else
"111111111111" when X = 272 AND Y = 99 else
"111111111111" when X = 273 AND Y = 99 else
"111111111111" when X = 274 AND Y = 99 else
"110111011111" when X = 275 AND Y = 99 else
"110111011111" when X = 276 AND Y = 99 else
"110111011111" when X = 277 AND Y = 99 else
"110111011111" when X = 278 AND Y = 99 else
"110111011111" when X = 279 AND Y = 99 else
"110111011111" when X = 280 AND Y = 99 else
"110111011111" when X = 281 AND Y = 99 else
"110111011111" when X = 282 AND Y = 99 else
"110111011111" when X = 283 AND Y = 99 else
"110111011111" when X = 284 AND Y = 99 else
"111111111111" when X = 285 AND Y = 99 else
"111111111111" when X = 286 AND Y = 99 else
"111111111111" when X = 287 AND Y = 99 else
"111111111111" when X = 288 AND Y = 99 else
"111111111111" when X = 289 AND Y = 99 else
"111111111111" when X = 290 AND Y = 99 else
"111111111111" when X = 291 AND Y = 99 else
"111111111111" when X = 292 AND Y = 99 else
"111111111111" when X = 293 AND Y = 99 else
"111111111111" when X = 294 AND Y = 99 else
"111111111111" when X = 295 AND Y = 99 else
"111111111111" when X = 296 AND Y = 99 else
"111111111111" when X = 297 AND Y = 99 else
"111111111111" when X = 298 AND Y = 99 else
"111111111111" when X = 299 AND Y = 99 else
"111111111111" when X = 300 AND Y = 99 else
"111111111111" when X = 301 AND Y = 99 else
"111111111111" when X = 302 AND Y = 99 else
"111111111111" when X = 303 AND Y = 99 else
"111111111111" when X = 304 AND Y = 99 else
"110111011111" when X = 305 AND Y = 99 else
"110111011111" when X = 306 AND Y = 99 else
"110111011111" when X = 307 AND Y = 99 else
"110111011111" when X = 308 AND Y = 99 else
"110111011111" when X = 309 AND Y = 99 else
"110111011111" when X = 310 AND Y = 99 else
"110111011111" when X = 311 AND Y = 99 else
"110111011111" when X = 312 AND Y = 99 else
"110111011111" when X = 313 AND Y = 99 else
"110111011111" when X = 314 AND Y = 99 else
"110111011111" when X = 315 AND Y = 99 else
"110111011111" when X = 316 AND Y = 99 else
"110111011111" when X = 317 AND Y = 99 else
"110111011111" when X = 318 AND Y = 99 else
"110111011111" when X = 319 AND Y = 99 else
"110111011111" when X = 320 AND Y = 99 else
"110111011111" when X = 321 AND Y = 99 else
"110111011111" when X = 322 AND Y = 99 else
"110111011111" when X = 323 AND Y = 99 else
"110111011111" when X = 324 AND Y = 99 else
"100010011101" when X = 0 AND Y = 100 else
"100010011101" when X = 1 AND Y = 100 else
"100010011101" when X = 2 AND Y = 100 else
"100010011101" when X = 3 AND Y = 100 else
"100010011101" when X = 4 AND Y = 100 else
"100010011101" when X = 5 AND Y = 100 else
"100010011101" when X = 6 AND Y = 100 else
"100010011101" when X = 7 AND Y = 100 else
"100010011101" when X = 8 AND Y = 100 else
"100010011101" when X = 9 AND Y = 100 else
"100010011101" when X = 10 AND Y = 100 else
"100010011101" when X = 11 AND Y = 100 else
"100010011101" when X = 12 AND Y = 100 else
"100010011101" when X = 13 AND Y = 100 else
"100010011101" when X = 14 AND Y = 100 else
"100010011101" when X = 15 AND Y = 100 else
"100010011101" when X = 16 AND Y = 100 else
"100010011101" when X = 17 AND Y = 100 else
"100010011101" when X = 18 AND Y = 100 else
"100010011101" when X = 19 AND Y = 100 else
"110111011111" when X = 20 AND Y = 100 else
"110111011111" when X = 21 AND Y = 100 else
"110111011111" when X = 22 AND Y = 100 else
"110111011111" when X = 23 AND Y = 100 else
"110111011111" when X = 24 AND Y = 100 else
"110111011111" when X = 25 AND Y = 100 else
"110111011111" when X = 26 AND Y = 100 else
"110111011111" when X = 27 AND Y = 100 else
"110111011111" when X = 28 AND Y = 100 else
"110111011111" when X = 29 AND Y = 100 else
"110111011111" when X = 30 AND Y = 100 else
"110111011111" when X = 31 AND Y = 100 else
"110111011111" when X = 32 AND Y = 100 else
"110111011111" when X = 33 AND Y = 100 else
"110111011111" when X = 34 AND Y = 100 else
"110111011111" when X = 35 AND Y = 100 else
"110111011111" when X = 36 AND Y = 100 else
"110111011111" when X = 37 AND Y = 100 else
"110111011111" when X = 38 AND Y = 100 else
"110111011111" when X = 39 AND Y = 100 else
"110111011111" when X = 40 AND Y = 100 else
"110111011111" when X = 41 AND Y = 100 else
"110111011111" when X = 42 AND Y = 100 else
"110111011111" when X = 43 AND Y = 100 else
"110111011111" when X = 44 AND Y = 100 else
"110111011111" when X = 45 AND Y = 100 else
"110111011111" when X = 46 AND Y = 100 else
"110111011111" when X = 47 AND Y = 100 else
"110111011111" when X = 48 AND Y = 100 else
"110111011111" when X = 49 AND Y = 100 else
"110111011111" when X = 50 AND Y = 100 else
"110111011111" when X = 51 AND Y = 100 else
"110111011111" when X = 52 AND Y = 100 else
"110111011111" when X = 53 AND Y = 100 else
"110111011111" when X = 54 AND Y = 100 else
"110111011111" when X = 55 AND Y = 100 else
"110111011111" when X = 56 AND Y = 100 else
"110111011111" when X = 57 AND Y = 100 else
"110111011111" when X = 58 AND Y = 100 else
"110111011111" when X = 59 AND Y = 100 else
"110111011111" when X = 60 AND Y = 100 else
"110111011111" when X = 61 AND Y = 100 else
"110111011111" when X = 62 AND Y = 100 else
"110111011111" when X = 63 AND Y = 100 else
"110111011111" when X = 64 AND Y = 100 else
"110111011111" when X = 65 AND Y = 100 else
"110111011111" when X = 66 AND Y = 100 else
"110111011111" when X = 67 AND Y = 100 else
"110111011111" when X = 68 AND Y = 100 else
"110111011111" when X = 69 AND Y = 100 else
"111111111111" when X = 70 AND Y = 100 else
"111111111111" when X = 71 AND Y = 100 else
"111111111111" when X = 72 AND Y = 100 else
"111111111111" when X = 73 AND Y = 100 else
"111111111111" when X = 74 AND Y = 100 else
"111111111111" when X = 75 AND Y = 100 else
"111111111111" when X = 76 AND Y = 100 else
"111111111111" when X = 77 AND Y = 100 else
"111111111111" when X = 78 AND Y = 100 else
"111111111111" when X = 79 AND Y = 100 else
"111111111111" when X = 80 AND Y = 100 else
"111111111111" when X = 81 AND Y = 100 else
"111111111111" when X = 82 AND Y = 100 else
"111111111111" when X = 83 AND Y = 100 else
"111111111111" when X = 84 AND Y = 100 else
"111111111111" when X = 85 AND Y = 100 else
"111111111111" when X = 86 AND Y = 100 else
"111111111111" when X = 87 AND Y = 100 else
"111111111111" when X = 88 AND Y = 100 else
"111111111111" when X = 89 AND Y = 100 else
"111111111111" when X = 90 AND Y = 100 else
"111111111111" when X = 91 AND Y = 100 else
"111111111111" when X = 92 AND Y = 100 else
"111111111111" when X = 93 AND Y = 100 else
"111111111111" when X = 94 AND Y = 100 else
"111111111111" when X = 95 AND Y = 100 else
"111111111111" when X = 96 AND Y = 100 else
"111111111111" when X = 97 AND Y = 100 else
"111111111111" when X = 98 AND Y = 100 else
"111111111111" when X = 99 AND Y = 100 else
"111111111111" when X = 100 AND Y = 100 else
"111111111111" when X = 101 AND Y = 100 else
"111111111111" when X = 102 AND Y = 100 else
"111111111111" when X = 103 AND Y = 100 else
"111111111111" when X = 104 AND Y = 100 else
"111111111111" when X = 105 AND Y = 100 else
"111111111111" when X = 106 AND Y = 100 else
"111111111111" when X = 107 AND Y = 100 else
"111111111111" when X = 108 AND Y = 100 else
"111111111111" when X = 109 AND Y = 100 else
"111111111111" when X = 110 AND Y = 100 else
"111111111111" when X = 111 AND Y = 100 else
"111111111111" when X = 112 AND Y = 100 else
"111111111111" when X = 113 AND Y = 100 else
"111111111111" when X = 114 AND Y = 100 else
"111111111111" when X = 115 AND Y = 100 else
"111111111111" when X = 116 AND Y = 100 else
"111111111111" when X = 117 AND Y = 100 else
"111111111111" when X = 118 AND Y = 100 else
"111111111111" when X = 119 AND Y = 100 else
"111111111111" when X = 120 AND Y = 100 else
"111111111111" when X = 121 AND Y = 100 else
"111111111111" when X = 122 AND Y = 100 else
"111111111111" when X = 123 AND Y = 100 else
"111111111111" when X = 124 AND Y = 100 else
"111111111111" when X = 125 AND Y = 100 else
"111111111111" when X = 126 AND Y = 100 else
"111111111111" when X = 127 AND Y = 100 else
"111111111111" when X = 128 AND Y = 100 else
"111111111111" when X = 129 AND Y = 100 else
"111111111111" when X = 130 AND Y = 100 else
"111111111111" when X = 131 AND Y = 100 else
"111111111111" when X = 132 AND Y = 100 else
"111111111111" when X = 133 AND Y = 100 else
"111111111111" when X = 134 AND Y = 100 else
"111111111111" when X = 135 AND Y = 100 else
"111111111111" when X = 136 AND Y = 100 else
"111111111111" when X = 137 AND Y = 100 else
"111111111111" when X = 138 AND Y = 100 else
"111111111111" when X = 139 AND Y = 100 else
"111111111111" when X = 140 AND Y = 100 else
"111111111111" when X = 141 AND Y = 100 else
"111111111111" when X = 142 AND Y = 100 else
"111111111111" when X = 143 AND Y = 100 else
"111111111111" when X = 144 AND Y = 100 else
"111111111111" when X = 145 AND Y = 100 else
"111111111111" when X = 146 AND Y = 100 else
"111111111111" when X = 147 AND Y = 100 else
"111111111111" when X = 148 AND Y = 100 else
"111111111111" when X = 149 AND Y = 100 else
"111111111111" when X = 150 AND Y = 100 else
"111111111111" when X = 151 AND Y = 100 else
"111111111111" when X = 152 AND Y = 100 else
"111111111111" when X = 153 AND Y = 100 else
"111111111111" when X = 154 AND Y = 100 else
"111111111111" when X = 155 AND Y = 100 else
"111111111111" when X = 156 AND Y = 100 else
"111111111111" when X = 157 AND Y = 100 else
"111111111111" when X = 158 AND Y = 100 else
"111111111111" when X = 159 AND Y = 100 else
"110111011111" when X = 160 AND Y = 100 else
"110111011111" when X = 161 AND Y = 100 else
"110111011111" when X = 162 AND Y = 100 else
"110111011111" when X = 163 AND Y = 100 else
"110111011111" when X = 164 AND Y = 100 else
"110111011111" when X = 165 AND Y = 100 else
"110111011111" when X = 166 AND Y = 100 else
"110111011111" when X = 167 AND Y = 100 else
"110111011111" when X = 168 AND Y = 100 else
"110111011111" when X = 169 AND Y = 100 else
"110111011111" when X = 170 AND Y = 100 else
"110111011111" when X = 171 AND Y = 100 else
"110111011111" when X = 172 AND Y = 100 else
"110111011111" when X = 173 AND Y = 100 else
"110111011111" when X = 174 AND Y = 100 else
"110111011111" when X = 175 AND Y = 100 else
"110111011111" when X = 176 AND Y = 100 else
"110111011111" when X = 177 AND Y = 100 else
"110111011111" when X = 178 AND Y = 100 else
"110111011111" when X = 179 AND Y = 100 else
"110111011111" when X = 180 AND Y = 100 else
"110111011111" when X = 181 AND Y = 100 else
"110111011111" when X = 182 AND Y = 100 else
"110111011111" when X = 183 AND Y = 100 else
"110111011111" when X = 184 AND Y = 100 else
"110111011111" when X = 185 AND Y = 100 else
"110111011111" when X = 186 AND Y = 100 else
"110111011111" when X = 187 AND Y = 100 else
"110111011111" when X = 188 AND Y = 100 else
"110111011111" when X = 189 AND Y = 100 else
"110111011111" when X = 190 AND Y = 100 else
"110111011111" when X = 191 AND Y = 100 else
"110111011111" when X = 192 AND Y = 100 else
"110111011111" when X = 193 AND Y = 100 else
"110111011111" when X = 194 AND Y = 100 else
"110111011111" when X = 195 AND Y = 100 else
"110111011111" when X = 196 AND Y = 100 else
"110111011111" when X = 197 AND Y = 100 else
"110111011111" when X = 198 AND Y = 100 else
"110111011111" when X = 199 AND Y = 100 else
"110111011111" when X = 200 AND Y = 100 else
"110111011111" when X = 201 AND Y = 100 else
"110111011111" when X = 202 AND Y = 100 else
"110111011111" when X = 203 AND Y = 100 else
"110111011111" when X = 204 AND Y = 100 else
"110111011111" when X = 205 AND Y = 100 else
"110111011111" when X = 206 AND Y = 100 else
"110111011111" when X = 207 AND Y = 100 else
"110111011111" when X = 208 AND Y = 100 else
"110111011111" when X = 209 AND Y = 100 else
"110111011111" when X = 210 AND Y = 100 else
"110111011111" when X = 211 AND Y = 100 else
"110111011111" when X = 212 AND Y = 100 else
"110111011111" when X = 213 AND Y = 100 else
"110111011111" when X = 214 AND Y = 100 else
"111111111111" when X = 215 AND Y = 100 else
"111111111111" when X = 216 AND Y = 100 else
"111111111111" when X = 217 AND Y = 100 else
"111111111111" when X = 218 AND Y = 100 else
"111111111111" when X = 219 AND Y = 100 else
"111111111111" when X = 220 AND Y = 100 else
"111111111111" when X = 221 AND Y = 100 else
"111111111111" when X = 222 AND Y = 100 else
"111111111111" when X = 223 AND Y = 100 else
"111111111111" when X = 224 AND Y = 100 else
"111111111111" when X = 225 AND Y = 100 else
"111111111111" when X = 226 AND Y = 100 else
"111111111111" when X = 227 AND Y = 100 else
"111111111111" when X = 228 AND Y = 100 else
"111111111111" when X = 229 AND Y = 100 else
"111111111111" when X = 230 AND Y = 100 else
"111111111111" when X = 231 AND Y = 100 else
"111111111111" when X = 232 AND Y = 100 else
"111111111111" when X = 233 AND Y = 100 else
"111111111111" when X = 234 AND Y = 100 else
"111111111111" when X = 235 AND Y = 100 else
"111111111111" when X = 236 AND Y = 100 else
"111111111111" when X = 237 AND Y = 100 else
"111111111111" when X = 238 AND Y = 100 else
"111111111111" when X = 239 AND Y = 100 else
"110111011111" when X = 240 AND Y = 100 else
"110111011111" when X = 241 AND Y = 100 else
"110111011111" when X = 242 AND Y = 100 else
"110111011111" when X = 243 AND Y = 100 else
"110111011111" when X = 244 AND Y = 100 else
"110111011111" when X = 245 AND Y = 100 else
"110111011111" when X = 246 AND Y = 100 else
"110111011111" when X = 247 AND Y = 100 else
"110111011111" when X = 248 AND Y = 100 else
"110111011111" when X = 249 AND Y = 100 else
"111111111111" when X = 250 AND Y = 100 else
"111111111111" when X = 251 AND Y = 100 else
"111111111111" when X = 252 AND Y = 100 else
"111111111111" when X = 253 AND Y = 100 else
"111111111111" when X = 254 AND Y = 100 else
"111111111111" when X = 255 AND Y = 100 else
"111111111111" when X = 256 AND Y = 100 else
"111111111111" when X = 257 AND Y = 100 else
"111111111111" when X = 258 AND Y = 100 else
"111111111111" when X = 259 AND Y = 100 else
"111111111111" when X = 260 AND Y = 100 else
"111111111111" when X = 261 AND Y = 100 else
"111111111111" when X = 262 AND Y = 100 else
"111111111111" when X = 263 AND Y = 100 else
"111111111111" when X = 264 AND Y = 100 else
"111111111111" when X = 265 AND Y = 100 else
"111111111111" when X = 266 AND Y = 100 else
"111111111111" when X = 267 AND Y = 100 else
"111111111111" when X = 268 AND Y = 100 else
"111111111111" when X = 269 AND Y = 100 else
"111111111111" when X = 270 AND Y = 100 else
"111111111111" when X = 271 AND Y = 100 else
"111111111111" when X = 272 AND Y = 100 else
"111111111111" when X = 273 AND Y = 100 else
"111111111111" when X = 274 AND Y = 100 else
"110111011111" when X = 275 AND Y = 100 else
"110111011111" when X = 276 AND Y = 100 else
"110111011111" when X = 277 AND Y = 100 else
"110111011111" when X = 278 AND Y = 100 else
"110111011111" when X = 279 AND Y = 100 else
"111111111111" when X = 280 AND Y = 100 else
"111111111111" when X = 281 AND Y = 100 else
"111111111111" when X = 282 AND Y = 100 else
"111111111111" when X = 283 AND Y = 100 else
"111111111111" when X = 284 AND Y = 100 else
"111111111111" when X = 285 AND Y = 100 else
"111111111111" when X = 286 AND Y = 100 else
"111111111111" when X = 287 AND Y = 100 else
"111111111111" when X = 288 AND Y = 100 else
"111111111111" when X = 289 AND Y = 100 else
"111111111111" when X = 290 AND Y = 100 else
"111111111111" when X = 291 AND Y = 100 else
"111111111111" when X = 292 AND Y = 100 else
"111111111111" when X = 293 AND Y = 100 else
"111111111111" when X = 294 AND Y = 100 else
"111111111111" when X = 295 AND Y = 100 else
"111111111111" when X = 296 AND Y = 100 else
"111111111111" when X = 297 AND Y = 100 else
"111111111111" when X = 298 AND Y = 100 else
"111111111111" when X = 299 AND Y = 100 else
"111111111111" when X = 300 AND Y = 100 else
"111111111111" when X = 301 AND Y = 100 else
"111111111111" when X = 302 AND Y = 100 else
"111111111111" when X = 303 AND Y = 100 else
"111111111111" when X = 304 AND Y = 100 else
"110111011111" when X = 305 AND Y = 100 else
"110111011111" when X = 306 AND Y = 100 else
"110111011111" when X = 307 AND Y = 100 else
"110111011111" when X = 308 AND Y = 100 else
"110111011111" when X = 309 AND Y = 100 else
"110111011111" when X = 310 AND Y = 100 else
"110111011111" when X = 311 AND Y = 100 else
"110111011111" when X = 312 AND Y = 100 else
"110111011111" when X = 313 AND Y = 100 else
"110111011111" when X = 314 AND Y = 100 else
"110111011111" when X = 315 AND Y = 100 else
"110111011111" when X = 316 AND Y = 100 else
"110111011111" when X = 317 AND Y = 100 else
"110111011111" when X = 318 AND Y = 100 else
"110111011111" when X = 319 AND Y = 100 else
"110111011111" when X = 320 AND Y = 100 else
"110111011111" when X = 321 AND Y = 100 else
"110111011111" when X = 322 AND Y = 100 else
"110111011111" when X = 323 AND Y = 100 else
"110111011111" when X = 324 AND Y = 100 else
"100010011101" when X = 0 AND Y = 101 else
"100010011101" when X = 1 AND Y = 101 else
"100010011101" when X = 2 AND Y = 101 else
"100010011101" when X = 3 AND Y = 101 else
"100010011101" when X = 4 AND Y = 101 else
"100010011101" when X = 5 AND Y = 101 else
"100010011101" when X = 6 AND Y = 101 else
"100010011101" when X = 7 AND Y = 101 else
"100010011101" when X = 8 AND Y = 101 else
"100010011101" when X = 9 AND Y = 101 else
"100010011101" when X = 10 AND Y = 101 else
"100010011101" when X = 11 AND Y = 101 else
"100010011101" when X = 12 AND Y = 101 else
"100010011101" when X = 13 AND Y = 101 else
"100010011101" when X = 14 AND Y = 101 else
"100010011101" when X = 15 AND Y = 101 else
"100010011101" when X = 16 AND Y = 101 else
"100010011101" when X = 17 AND Y = 101 else
"100010011101" when X = 18 AND Y = 101 else
"100010011101" when X = 19 AND Y = 101 else
"110111011111" when X = 20 AND Y = 101 else
"110111011111" when X = 21 AND Y = 101 else
"110111011111" when X = 22 AND Y = 101 else
"110111011111" when X = 23 AND Y = 101 else
"110111011111" when X = 24 AND Y = 101 else
"110111011111" when X = 25 AND Y = 101 else
"110111011111" when X = 26 AND Y = 101 else
"110111011111" when X = 27 AND Y = 101 else
"110111011111" when X = 28 AND Y = 101 else
"110111011111" when X = 29 AND Y = 101 else
"110111011111" when X = 30 AND Y = 101 else
"110111011111" when X = 31 AND Y = 101 else
"110111011111" when X = 32 AND Y = 101 else
"110111011111" when X = 33 AND Y = 101 else
"110111011111" when X = 34 AND Y = 101 else
"110111011111" when X = 35 AND Y = 101 else
"110111011111" when X = 36 AND Y = 101 else
"110111011111" when X = 37 AND Y = 101 else
"110111011111" when X = 38 AND Y = 101 else
"110111011111" when X = 39 AND Y = 101 else
"110111011111" when X = 40 AND Y = 101 else
"110111011111" when X = 41 AND Y = 101 else
"110111011111" when X = 42 AND Y = 101 else
"110111011111" when X = 43 AND Y = 101 else
"110111011111" when X = 44 AND Y = 101 else
"110111011111" when X = 45 AND Y = 101 else
"110111011111" when X = 46 AND Y = 101 else
"110111011111" when X = 47 AND Y = 101 else
"110111011111" when X = 48 AND Y = 101 else
"110111011111" when X = 49 AND Y = 101 else
"110111011111" when X = 50 AND Y = 101 else
"110111011111" when X = 51 AND Y = 101 else
"110111011111" when X = 52 AND Y = 101 else
"110111011111" when X = 53 AND Y = 101 else
"110111011111" when X = 54 AND Y = 101 else
"110111011111" when X = 55 AND Y = 101 else
"110111011111" when X = 56 AND Y = 101 else
"110111011111" when X = 57 AND Y = 101 else
"110111011111" when X = 58 AND Y = 101 else
"110111011111" when X = 59 AND Y = 101 else
"110111011111" when X = 60 AND Y = 101 else
"110111011111" when X = 61 AND Y = 101 else
"110111011111" when X = 62 AND Y = 101 else
"110111011111" when X = 63 AND Y = 101 else
"110111011111" when X = 64 AND Y = 101 else
"110111011111" when X = 65 AND Y = 101 else
"110111011111" when X = 66 AND Y = 101 else
"110111011111" when X = 67 AND Y = 101 else
"110111011111" when X = 68 AND Y = 101 else
"110111011111" when X = 69 AND Y = 101 else
"111111111111" when X = 70 AND Y = 101 else
"111111111111" when X = 71 AND Y = 101 else
"111111111111" when X = 72 AND Y = 101 else
"111111111111" when X = 73 AND Y = 101 else
"111111111111" when X = 74 AND Y = 101 else
"111111111111" when X = 75 AND Y = 101 else
"111111111111" when X = 76 AND Y = 101 else
"111111111111" when X = 77 AND Y = 101 else
"111111111111" when X = 78 AND Y = 101 else
"111111111111" when X = 79 AND Y = 101 else
"111111111111" when X = 80 AND Y = 101 else
"111111111111" when X = 81 AND Y = 101 else
"111111111111" when X = 82 AND Y = 101 else
"111111111111" when X = 83 AND Y = 101 else
"111111111111" when X = 84 AND Y = 101 else
"111111111111" when X = 85 AND Y = 101 else
"111111111111" when X = 86 AND Y = 101 else
"111111111111" when X = 87 AND Y = 101 else
"111111111111" when X = 88 AND Y = 101 else
"111111111111" when X = 89 AND Y = 101 else
"111111111111" when X = 90 AND Y = 101 else
"111111111111" when X = 91 AND Y = 101 else
"111111111111" when X = 92 AND Y = 101 else
"111111111111" when X = 93 AND Y = 101 else
"111111111111" when X = 94 AND Y = 101 else
"111111111111" when X = 95 AND Y = 101 else
"111111111111" when X = 96 AND Y = 101 else
"111111111111" when X = 97 AND Y = 101 else
"111111111111" when X = 98 AND Y = 101 else
"111111111111" when X = 99 AND Y = 101 else
"111111111111" when X = 100 AND Y = 101 else
"111111111111" when X = 101 AND Y = 101 else
"111111111111" when X = 102 AND Y = 101 else
"111111111111" when X = 103 AND Y = 101 else
"111111111111" when X = 104 AND Y = 101 else
"111111111111" when X = 105 AND Y = 101 else
"111111111111" when X = 106 AND Y = 101 else
"111111111111" when X = 107 AND Y = 101 else
"111111111111" when X = 108 AND Y = 101 else
"111111111111" when X = 109 AND Y = 101 else
"111111111111" when X = 110 AND Y = 101 else
"111111111111" when X = 111 AND Y = 101 else
"111111111111" when X = 112 AND Y = 101 else
"111111111111" when X = 113 AND Y = 101 else
"111111111111" when X = 114 AND Y = 101 else
"111111111111" when X = 115 AND Y = 101 else
"111111111111" when X = 116 AND Y = 101 else
"111111111111" when X = 117 AND Y = 101 else
"111111111111" when X = 118 AND Y = 101 else
"111111111111" when X = 119 AND Y = 101 else
"111111111111" when X = 120 AND Y = 101 else
"111111111111" when X = 121 AND Y = 101 else
"111111111111" when X = 122 AND Y = 101 else
"111111111111" when X = 123 AND Y = 101 else
"111111111111" when X = 124 AND Y = 101 else
"111111111111" when X = 125 AND Y = 101 else
"111111111111" when X = 126 AND Y = 101 else
"111111111111" when X = 127 AND Y = 101 else
"111111111111" when X = 128 AND Y = 101 else
"111111111111" when X = 129 AND Y = 101 else
"111111111111" when X = 130 AND Y = 101 else
"111111111111" when X = 131 AND Y = 101 else
"111111111111" when X = 132 AND Y = 101 else
"111111111111" when X = 133 AND Y = 101 else
"111111111111" when X = 134 AND Y = 101 else
"111111111111" when X = 135 AND Y = 101 else
"111111111111" when X = 136 AND Y = 101 else
"111111111111" when X = 137 AND Y = 101 else
"111111111111" when X = 138 AND Y = 101 else
"111111111111" when X = 139 AND Y = 101 else
"111111111111" when X = 140 AND Y = 101 else
"111111111111" when X = 141 AND Y = 101 else
"111111111111" when X = 142 AND Y = 101 else
"111111111111" when X = 143 AND Y = 101 else
"111111111111" when X = 144 AND Y = 101 else
"111111111111" when X = 145 AND Y = 101 else
"111111111111" when X = 146 AND Y = 101 else
"111111111111" when X = 147 AND Y = 101 else
"111111111111" when X = 148 AND Y = 101 else
"111111111111" when X = 149 AND Y = 101 else
"111111111111" when X = 150 AND Y = 101 else
"111111111111" when X = 151 AND Y = 101 else
"111111111111" when X = 152 AND Y = 101 else
"111111111111" when X = 153 AND Y = 101 else
"111111111111" when X = 154 AND Y = 101 else
"111111111111" when X = 155 AND Y = 101 else
"111111111111" when X = 156 AND Y = 101 else
"111111111111" when X = 157 AND Y = 101 else
"111111111111" when X = 158 AND Y = 101 else
"111111111111" when X = 159 AND Y = 101 else
"110111011111" when X = 160 AND Y = 101 else
"110111011111" when X = 161 AND Y = 101 else
"110111011111" when X = 162 AND Y = 101 else
"110111011111" when X = 163 AND Y = 101 else
"110111011111" when X = 164 AND Y = 101 else
"110111011111" when X = 165 AND Y = 101 else
"110111011111" when X = 166 AND Y = 101 else
"110111011111" when X = 167 AND Y = 101 else
"110111011111" when X = 168 AND Y = 101 else
"110111011111" when X = 169 AND Y = 101 else
"110111011111" when X = 170 AND Y = 101 else
"110111011111" when X = 171 AND Y = 101 else
"110111011111" when X = 172 AND Y = 101 else
"110111011111" when X = 173 AND Y = 101 else
"110111011111" when X = 174 AND Y = 101 else
"110111011111" when X = 175 AND Y = 101 else
"110111011111" when X = 176 AND Y = 101 else
"110111011111" when X = 177 AND Y = 101 else
"110111011111" when X = 178 AND Y = 101 else
"110111011111" when X = 179 AND Y = 101 else
"110111011111" when X = 180 AND Y = 101 else
"110111011111" when X = 181 AND Y = 101 else
"110111011111" when X = 182 AND Y = 101 else
"110111011111" when X = 183 AND Y = 101 else
"110111011111" when X = 184 AND Y = 101 else
"110111011111" when X = 185 AND Y = 101 else
"110111011111" when X = 186 AND Y = 101 else
"110111011111" when X = 187 AND Y = 101 else
"110111011111" when X = 188 AND Y = 101 else
"110111011111" when X = 189 AND Y = 101 else
"110111011111" when X = 190 AND Y = 101 else
"110111011111" when X = 191 AND Y = 101 else
"110111011111" when X = 192 AND Y = 101 else
"110111011111" when X = 193 AND Y = 101 else
"110111011111" when X = 194 AND Y = 101 else
"110111011111" when X = 195 AND Y = 101 else
"110111011111" when X = 196 AND Y = 101 else
"110111011111" when X = 197 AND Y = 101 else
"110111011111" when X = 198 AND Y = 101 else
"110111011111" when X = 199 AND Y = 101 else
"110111011111" when X = 200 AND Y = 101 else
"110111011111" when X = 201 AND Y = 101 else
"110111011111" when X = 202 AND Y = 101 else
"110111011111" when X = 203 AND Y = 101 else
"110111011111" when X = 204 AND Y = 101 else
"110111011111" when X = 205 AND Y = 101 else
"110111011111" when X = 206 AND Y = 101 else
"110111011111" when X = 207 AND Y = 101 else
"110111011111" when X = 208 AND Y = 101 else
"110111011111" when X = 209 AND Y = 101 else
"110111011111" when X = 210 AND Y = 101 else
"110111011111" when X = 211 AND Y = 101 else
"110111011111" when X = 212 AND Y = 101 else
"110111011111" when X = 213 AND Y = 101 else
"110111011111" when X = 214 AND Y = 101 else
"111111111111" when X = 215 AND Y = 101 else
"111111111111" when X = 216 AND Y = 101 else
"111111111111" when X = 217 AND Y = 101 else
"111111111111" when X = 218 AND Y = 101 else
"111111111111" when X = 219 AND Y = 101 else
"111111111111" when X = 220 AND Y = 101 else
"111111111111" when X = 221 AND Y = 101 else
"111111111111" when X = 222 AND Y = 101 else
"111111111111" when X = 223 AND Y = 101 else
"111111111111" when X = 224 AND Y = 101 else
"111111111111" when X = 225 AND Y = 101 else
"111111111111" when X = 226 AND Y = 101 else
"111111111111" when X = 227 AND Y = 101 else
"111111111111" when X = 228 AND Y = 101 else
"111111111111" when X = 229 AND Y = 101 else
"111111111111" when X = 230 AND Y = 101 else
"111111111111" when X = 231 AND Y = 101 else
"111111111111" when X = 232 AND Y = 101 else
"111111111111" when X = 233 AND Y = 101 else
"111111111111" when X = 234 AND Y = 101 else
"111111111111" when X = 235 AND Y = 101 else
"111111111111" when X = 236 AND Y = 101 else
"111111111111" when X = 237 AND Y = 101 else
"111111111111" when X = 238 AND Y = 101 else
"111111111111" when X = 239 AND Y = 101 else
"110111011111" when X = 240 AND Y = 101 else
"110111011111" when X = 241 AND Y = 101 else
"110111011111" when X = 242 AND Y = 101 else
"110111011111" when X = 243 AND Y = 101 else
"110111011111" when X = 244 AND Y = 101 else
"110111011111" when X = 245 AND Y = 101 else
"110111011111" when X = 246 AND Y = 101 else
"110111011111" when X = 247 AND Y = 101 else
"110111011111" when X = 248 AND Y = 101 else
"110111011111" when X = 249 AND Y = 101 else
"111111111111" when X = 250 AND Y = 101 else
"111111111111" when X = 251 AND Y = 101 else
"111111111111" when X = 252 AND Y = 101 else
"111111111111" when X = 253 AND Y = 101 else
"111111111111" when X = 254 AND Y = 101 else
"111111111111" when X = 255 AND Y = 101 else
"111111111111" when X = 256 AND Y = 101 else
"111111111111" when X = 257 AND Y = 101 else
"111111111111" when X = 258 AND Y = 101 else
"111111111111" when X = 259 AND Y = 101 else
"111111111111" when X = 260 AND Y = 101 else
"111111111111" when X = 261 AND Y = 101 else
"111111111111" when X = 262 AND Y = 101 else
"111111111111" when X = 263 AND Y = 101 else
"111111111111" when X = 264 AND Y = 101 else
"111111111111" when X = 265 AND Y = 101 else
"111111111111" when X = 266 AND Y = 101 else
"111111111111" when X = 267 AND Y = 101 else
"111111111111" when X = 268 AND Y = 101 else
"111111111111" when X = 269 AND Y = 101 else
"111111111111" when X = 270 AND Y = 101 else
"111111111111" when X = 271 AND Y = 101 else
"111111111111" when X = 272 AND Y = 101 else
"111111111111" when X = 273 AND Y = 101 else
"111111111111" when X = 274 AND Y = 101 else
"110111011111" when X = 275 AND Y = 101 else
"110111011111" when X = 276 AND Y = 101 else
"110111011111" when X = 277 AND Y = 101 else
"110111011111" when X = 278 AND Y = 101 else
"110111011111" when X = 279 AND Y = 101 else
"111111111111" when X = 280 AND Y = 101 else
"111111111111" when X = 281 AND Y = 101 else
"111111111111" when X = 282 AND Y = 101 else
"111111111111" when X = 283 AND Y = 101 else
"111111111111" when X = 284 AND Y = 101 else
"111111111111" when X = 285 AND Y = 101 else
"111111111111" when X = 286 AND Y = 101 else
"111111111111" when X = 287 AND Y = 101 else
"111111111111" when X = 288 AND Y = 101 else
"111111111111" when X = 289 AND Y = 101 else
"111111111111" when X = 290 AND Y = 101 else
"111111111111" when X = 291 AND Y = 101 else
"111111111111" when X = 292 AND Y = 101 else
"111111111111" when X = 293 AND Y = 101 else
"111111111111" when X = 294 AND Y = 101 else
"111111111111" when X = 295 AND Y = 101 else
"111111111111" when X = 296 AND Y = 101 else
"111111111111" when X = 297 AND Y = 101 else
"111111111111" when X = 298 AND Y = 101 else
"111111111111" when X = 299 AND Y = 101 else
"111111111111" when X = 300 AND Y = 101 else
"111111111111" when X = 301 AND Y = 101 else
"111111111111" when X = 302 AND Y = 101 else
"111111111111" when X = 303 AND Y = 101 else
"111111111111" when X = 304 AND Y = 101 else
"110111011111" when X = 305 AND Y = 101 else
"110111011111" when X = 306 AND Y = 101 else
"110111011111" when X = 307 AND Y = 101 else
"110111011111" when X = 308 AND Y = 101 else
"110111011111" when X = 309 AND Y = 101 else
"110111011111" when X = 310 AND Y = 101 else
"110111011111" when X = 311 AND Y = 101 else
"110111011111" when X = 312 AND Y = 101 else
"110111011111" when X = 313 AND Y = 101 else
"110111011111" when X = 314 AND Y = 101 else
"110111011111" when X = 315 AND Y = 101 else
"110111011111" when X = 316 AND Y = 101 else
"110111011111" when X = 317 AND Y = 101 else
"110111011111" when X = 318 AND Y = 101 else
"110111011111" when X = 319 AND Y = 101 else
"110111011111" when X = 320 AND Y = 101 else
"110111011111" when X = 321 AND Y = 101 else
"110111011111" when X = 322 AND Y = 101 else
"110111011111" when X = 323 AND Y = 101 else
"110111011111" when X = 324 AND Y = 101 else
"100010011101" when X = 0 AND Y = 102 else
"100010011101" when X = 1 AND Y = 102 else
"100010011101" when X = 2 AND Y = 102 else
"100010011101" when X = 3 AND Y = 102 else
"100010011101" when X = 4 AND Y = 102 else
"100010011101" when X = 5 AND Y = 102 else
"100010011101" when X = 6 AND Y = 102 else
"100010011101" when X = 7 AND Y = 102 else
"100010011101" when X = 8 AND Y = 102 else
"100010011101" when X = 9 AND Y = 102 else
"100010011101" when X = 10 AND Y = 102 else
"100010011101" when X = 11 AND Y = 102 else
"100010011101" when X = 12 AND Y = 102 else
"100010011101" when X = 13 AND Y = 102 else
"100010011101" when X = 14 AND Y = 102 else
"100010011101" when X = 15 AND Y = 102 else
"100010011101" when X = 16 AND Y = 102 else
"100010011101" when X = 17 AND Y = 102 else
"100010011101" when X = 18 AND Y = 102 else
"100010011101" when X = 19 AND Y = 102 else
"110111011111" when X = 20 AND Y = 102 else
"110111011111" when X = 21 AND Y = 102 else
"110111011111" when X = 22 AND Y = 102 else
"110111011111" when X = 23 AND Y = 102 else
"110111011111" when X = 24 AND Y = 102 else
"110111011111" when X = 25 AND Y = 102 else
"110111011111" when X = 26 AND Y = 102 else
"110111011111" when X = 27 AND Y = 102 else
"110111011111" when X = 28 AND Y = 102 else
"110111011111" when X = 29 AND Y = 102 else
"110111011111" when X = 30 AND Y = 102 else
"110111011111" when X = 31 AND Y = 102 else
"110111011111" when X = 32 AND Y = 102 else
"110111011111" when X = 33 AND Y = 102 else
"110111011111" when X = 34 AND Y = 102 else
"110111011111" when X = 35 AND Y = 102 else
"110111011111" when X = 36 AND Y = 102 else
"110111011111" when X = 37 AND Y = 102 else
"110111011111" when X = 38 AND Y = 102 else
"110111011111" when X = 39 AND Y = 102 else
"110111011111" when X = 40 AND Y = 102 else
"110111011111" when X = 41 AND Y = 102 else
"110111011111" when X = 42 AND Y = 102 else
"110111011111" when X = 43 AND Y = 102 else
"110111011111" when X = 44 AND Y = 102 else
"110111011111" when X = 45 AND Y = 102 else
"110111011111" when X = 46 AND Y = 102 else
"110111011111" when X = 47 AND Y = 102 else
"110111011111" when X = 48 AND Y = 102 else
"110111011111" when X = 49 AND Y = 102 else
"110111011111" when X = 50 AND Y = 102 else
"110111011111" when X = 51 AND Y = 102 else
"110111011111" when X = 52 AND Y = 102 else
"110111011111" when X = 53 AND Y = 102 else
"110111011111" when X = 54 AND Y = 102 else
"110111011111" when X = 55 AND Y = 102 else
"110111011111" when X = 56 AND Y = 102 else
"110111011111" when X = 57 AND Y = 102 else
"110111011111" when X = 58 AND Y = 102 else
"110111011111" when X = 59 AND Y = 102 else
"110111011111" when X = 60 AND Y = 102 else
"110111011111" when X = 61 AND Y = 102 else
"110111011111" when X = 62 AND Y = 102 else
"110111011111" when X = 63 AND Y = 102 else
"110111011111" when X = 64 AND Y = 102 else
"110111011111" when X = 65 AND Y = 102 else
"110111011111" when X = 66 AND Y = 102 else
"110111011111" when X = 67 AND Y = 102 else
"110111011111" when X = 68 AND Y = 102 else
"110111011111" when X = 69 AND Y = 102 else
"111111111111" when X = 70 AND Y = 102 else
"111111111111" when X = 71 AND Y = 102 else
"111111111111" when X = 72 AND Y = 102 else
"111111111111" when X = 73 AND Y = 102 else
"111111111111" when X = 74 AND Y = 102 else
"111111111111" when X = 75 AND Y = 102 else
"111111111111" when X = 76 AND Y = 102 else
"111111111111" when X = 77 AND Y = 102 else
"111111111111" when X = 78 AND Y = 102 else
"111111111111" when X = 79 AND Y = 102 else
"111111111111" when X = 80 AND Y = 102 else
"111111111111" when X = 81 AND Y = 102 else
"111111111111" when X = 82 AND Y = 102 else
"111111111111" when X = 83 AND Y = 102 else
"111111111111" when X = 84 AND Y = 102 else
"111111111111" when X = 85 AND Y = 102 else
"111111111111" when X = 86 AND Y = 102 else
"111111111111" when X = 87 AND Y = 102 else
"111111111111" when X = 88 AND Y = 102 else
"111111111111" when X = 89 AND Y = 102 else
"111111111111" when X = 90 AND Y = 102 else
"111111111111" when X = 91 AND Y = 102 else
"111111111111" when X = 92 AND Y = 102 else
"111111111111" when X = 93 AND Y = 102 else
"111111111111" when X = 94 AND Y = 102 else
"111111111111" when X = 95 AND Y = 102 else
"111111111111" when X = 96 AND Y = 102 else
"111111111111" when X = 97 AND Y = 102 else
"111111111111" when X = 98 AND Y = 102 else
"111111111111" when X = 99 AND Y = 102 else
"111111111111" when X = 100 AND Y = 102 else
"111111111111" when X = 101 AND Y = 102 else
"111111111111" when X = 102 AND Y = 102 else
"111111111111" when X = 103 AND Y = 102 else
"111111111111" when X = 104 AND Y = 102 else
"111111111111" when X = 105 AND Y = 102 else
"111111111111" when X = 106 AND Y = 102 else
"111111111111" when X = 107 AND Y = 102 else
"111111111111" when X = 108 AND Y = 102 else
"111111111111" when X = 109 AND Y = 102 else
"111111111111" when X = 110 AND Y = 102 else
"111111111111" when X = 111 AND Y = 102 else
"111111111111" when X = 112 AND Y = 102 else
"111111111111" when X = 113 AND Y = 102 else
"111111111111" when X = 114 AND Y = 102 else
"111111111111" when X = 115 AND Y = 102 else
"111111111111" when X = 116 AND Y = 102 else
"111111111111" when X = 117 AND Y = 102 else
"111111111111" when X = 118 AND Y = 102 else
"111111111111" when X = 119 AND Y = 102 else
"111111111111" when X = 120 AND Y = 102 else
"111111111111" when X = 121 AND Y = 102 else
"111111111111" when X = 122 AND Y = 102 else
"111111111111" when X = 123 AND Y = 102 else
"111111111111" when X = 124 AND Y = 102 else
"111111111111" when X = 125 AND Y = 102 else
"111111111111" when X = 126 AND Y = 102 else
"111111111111" when X = 127 AND Y = 102 else
"111111111111" when X = 128 AND Y = 102 else
"111111111111" when X = 129 AND Y = 102 else
"111111111111" when X = 130 AND Y = 102 else
"111111111111" when X = 131 AND Y = 102 else
"111111111111" when X = 132 AND Y = 102 else
"111111111111" when X = 133 AND Y = 102 else
"111111111111" when X = 134 AND Y = 102 else
"111111111111" when X = 135 AND Y = 102 else
"111111111111" when X = 136 AND Y = 102 else
"111111111111" when X = 137 AND Y = 102 else
"111111111111" when X = 138 AND Y = 102 else
"111111111111" when X = 139 AND Y = 102 else
"111111111111" when X = 140 AND Y = 102 else
"111111111111" when X = 141 AND Y = 102 else
"111111111111" when X = 142 AND Y = 102 else
"111111111111" when X = 143 AND Y = 102 else
"111111111111" when X = 144 AND Y = 102 else
"111111111111" when X = 145 AND Y = 102 else
"111111111111" when X = 146 AND Y = 102 else
"111111111111" when X = 147 AND Y = 102 else
"111111111111" when X = 148 AND Y = 102 else
"111111111111" when X = 149 AND Y = 102 else
"111111111111" when X = 150 AND Y = 102 else
"111111111111" when X = 151 AND Y = 102 else
"111111111111" when X = 152 AND Y = 102 else
"111111111111" when X = 153 AND Y = 102 else
"111111111111" when X = 154 AND Y = 102 else
"111111111111" when X = 155 AND Y = 102 else
"111111111111" when X = 156 AND Y = 102 else
"111111111111" when X = 157 AND Y = 102 else
"111111111111" when X = 158 AND Y = 102 else
"111111111111" when X = 159 AND Y = 102 else
"110111011111" when X = 160 AND Y = 102 else
"110111011111" when X = 161 AND Y = 102 else
"110111011111" when X = 162 AND Y = 102 else
"110111011111" when X = 163 AND Y = 102 else
"110111011111" when X = 164 AND Y = 102 else
"110111011111" when X = 165 AND Y = 102 else
"110111011111" when X = 166 AND Y = 102 else
"110111011111" when X = 167 AND Y = 102 else
"110111011111" when X = 168 AND Y = 102 else
"110111011111" when X = 169 AND Y = 102 else
"110111011111" when X = 170 AND Y = 102 else
"110111011111" when X = 171 AND Y = 102 else
"110111011111" when X = 172 AND Y = 102 else
"110111011111" when X = 173 AND Y = 102 else
"110111011111" when X = 174 AND Y = 102 else
"110111011111" when X = 175 AND Y = 102 else
"110111011111" when X = 176 AND Y = 102 else
"110111011111" when X = 177 AND Y = 102 else
"110111011111" when X = 178 AND Y = 102 else
"110111011111" when X = 179 AND Y = 102 else
"110111011111" when X = 180 AND Y = 102 else
"110111011111" when X = 181 AND Y = 102 else
"110111011111" when X = 182 AND Y = 102 else
"110111011111" when X = 183 AND Y = 102 else
"110111011111" when X = 184 AND Y = 102 else
"110111011111" when X = 185 AND Y = 102 else
"110111011111" when X = 186 AND Y = 102 else
"110111011111" when X = 187 AND Y = 102 else
"110111011111" when X = 188 AND Y = 102 else
"110111011111" when X = 189 AND Y = 102 else
"110111011111" when X = 190 AND Y = 102 else
"110111011111" when X = 191 AND Y = 102 else
"110111011111" when X = 192 AND Y = 102 else
"110111011111" when X = 193 AND Y = 102 else
"110111011111" when X = 194 AND Y = 102 else
"110111011111" when X = 195 AND Y = 102 else
"110111011111" when X = 196 AND Y = 102 else
"110111011111" when X = 197 AND Y = 102 else
"110111011111" when X = 198 AND Y = 102 else
"110111011111" when X = 199 AND Y = 102 else
"110111011111" when X = 200 AND Y = 102 else
"110111011111" when X = 201 AND Y = 102 else
"110111011111" when X = 202 AND Y = 102 else
"110111011111" when X = 203 AND Y = 102 else
"110111011111" when X = 204 AND Y = 102 else
"110111011111" when X = 205 AND Y = 102 else
"110111011111" when X = 206 AND Y = 102 else
"110111011111" when X = 207 AND Y = 102 else
"110111011111" when X = 208 AND Y = 102 else
"110111011111" when X = 209 AND Y = 102 else
"110111011111" when X = 210 AND Y = 102 else
"110111011111" when X = 211 AND Y = 102 else
"110111011111" when X = 212 AND Y = 102 else
"110111011111" when X = 213 AND Y = 102 else
"110111011111" when X = 214 AND Y = 102 else
"111111111111" when X = 215 AND Y = 102 else
"111111111111" when X = 216 AND Y = 102 else
"111111111111" when X = 217 AND Y = 102 else
"111111111111" when X = 218 AND Y = 102 else
"111111111111" when X = 219 AND Y = 102 else
"111111111111" when X = 220 AND Y = 102 else
"111111111111" when X = 221 AND Y = 102 else
"111111111111" when X = 222 AND Y = 102 else
"111111111111" when X = 223 AND Y = 102 else
"111111111111" when X = 224 AND Y = 102 else
"111111111111" when X = 225 AND Y = 102 else
"111111111111" when X = 226 AND Y = 102 else
"111111111111" when X = 227 AND Y = 102 else
"111111111111" when X = 228 AND Y = 102 else
"111111111111" when X = 229 AND Y = 102 else
"111111111111" when X = 230 AND Y = 102 else
"111111111111" when X = 231 AND Y = 102 else
"111111111111" when X = 232 AND Y = 102 else
"111111111111" when X = 233 AND Y = 102 else
"111111111111" when X = 234 AND Y = 102 else
"111111111111" when X = 235 AND Y = 102 else
"111111111111" when X = 236 AND Y = 102 else
"111111111111" when X = 237 AND Y = 102 else
"111111111111" when X = 238 AND Y = 102 else
"111111111111" when X = 239 AND Y = 102 else
"110111011111" when X = 240 AND Y = 102 else
"110111011111" when X = 241 AND Y = 102 else
"110111011111" when X = 242 AND Y = 102 else
"110111011111" when X = 243 AND Y = 102 else
"110111011111" when X = 244 AND Y = 102 else
"110111011111" when X = 245 AND Y = 102 else
"110111011111" when X = 246 AND Y = 102 else
"110111011111" when X = 247 AND Y = 102 else
"110111011111" when X = 248 AND Y = 102 else
"110111011111" when X = 249 AND Y = 102 else
"111111111111" when X = 250 AND Y = 102 else
"111111111111" when X = 251 AND Y = 102 else
"111111111111" when X = 252 AND Y = 102 else
"111111111111" when X = 253 AND Y = 102 else
"111111111111" when X = 254 AND Y = 102 else
"111111111111" when X = 255 AND Y = 102 else
"111111111111" when X = 256 AND Y = 102 else
"111111111111" when X = 257 AND Y = 102 else
"111111111111" when X = 258 AND Y = 102 else
"111111111111" when X = 259 AND Y = 102 else
"111111111111" when X = 260 AND Y = 102 else
"111111111111" when X = 261 AND Y = 102 else
"111111111111" when X = 262 AND Y = 102 else
"111111111111" when X = 263 AND Y = 102 else
"111111111111" when X = 264 AND Y = 102 else
"111111111111" when X = 265 AND Y = 102 else
"111111111111" when X = 266 AND Y = 102 else
"111111111111" when X = 267 AND Y = 102 else
"111111111111" when X = 268 AND Y = 102 else
"111111111111" when X = 269 AND Y = 102 else
"111111111111" when X = 270 AND Y = 102 else
"111111111111" when X = 271 AND Y = 102 else
"111111111111" when X = 272 AND Y = 102 else
"111111111111" when X = 273 AND Y = 102 else
"111111111111" when X = 274 AND Y = 102 else
"110111011111" when X = 275 AND Y = 102 else
"110111011111" when X = 276 AND Y = 102 else
"110111011111" when X = 277 AND Y = 102 else
"110111011111" when X = 278 AND Y = 102 else
"110111011111" when X = 279 AND Y = 102 else
"111111111111" when X = 280 AND Y = 102 else
"111111111111" when X = 281 AND Y = 102 else
"111111111111" when X = 282 AND Y = 102 else
"111111111111" when X = 283 AND Y = 102 else
"111111111111" when X = 284 AND Y = 102 else
"111111111111" when X = 285 AND Y = 102 else
"111111111111" when X = 286 AND Y = 102 else
"111111111111" when X = 287 AND Y = 102 else
"111111111111" when X = 288 AND Y = 102 else
"111111111111" when X = 289 AND Y = 102 else
"111111111111" when X = 290 AND Y = 102 else
"111111111111" when X = 291 AND Y = 102 else
"111111111111" when X = 292 AND Y = 102 else
"111111111111" when X = 293 AND Y = 102 else
"111111111111" when X = 294 AND Y = 102 else
"111111111111" when X = 295 AND Y = 102 else
"111111111111" when X = 296 AND Y = 102 else
"111111111111" when X = 297 AND Y = 102 else
"111111111111" when X = 298 AND Y = 102 else
"111111111111" when X = 299 AND Y = 102 else
"111111111111" when X = 300 AND Y = 102 else
"111111111111" when X = 301 AND Y = 102 else
"111111111111" when X = 302 AND Y = 102 else
"111111111111" when X = 303 AND Y = 102 else
"111111111111" when X = 304 AND Y = 102 else
"110111011111" when X = 305 AND Y = 102 else
"110111011111" when X = 306 AND Y = 102 else
"110111011111" when X = 307 AND Y = 102 else
"110111011111" when X = 308 AND Y = 102 else
"110111011111" when X = 309 AND Y = 102 else
"110111011111" when X = 310 AND Y = 102 else
"110111011111" when X = 311 AND Y = 102 else
"110111011111" when X = 312 AND Y = 102 else
"110111011111" when X = 313 AND Y = 102 else
"110111011111" when X = 314 AND Y = 102 else
"110111011111" when X = 315 AND Y = 102 else
"110111011111" when X = 316 AND Y = 102 else
"110111011111" when X = 317 AND Y = 102 else
"110111011111" when X = 318 AND Y = 102 else
"110111011111" when X = 319 AND Y = 102 else
"110111011111" when X = 320 AND Y = 102 else
"110111011111" when X = 321 AND Y = 102 else
"110111011111" when X = 322 AND Y = 102 else
"110111011111" when X = 323 AND Y = 102 else
"110111011111" when X = 324 AND Y = 102 else
"100010011101" when X = 0 AND Y = 103 else
"100010011101" when X = 1 AND Y = 103 else
"100010011101" when X = 2 AND Y = 103 else
"100010011101" when X = 3 AND Y = 103 else
"100010011101" when X = 4 AND Y = 103 else
"100010011101" when X = 5 AND Y = 103 else
"100010011101" when X = 6 AND Y = 103 else
"100010011101" when X = 7 AND Y = 103 else
"100010011101" when X = 8 AND Y = 103 else
"100010011101" when X = 9 AND Y = 103 else
"100010011101" when X = 10 AND Y = 103 else
"100010011101" when X = 11 AND Y = 103 else
"100010011101" when X = 12 AND Y = 103 else
"100010011101" when X = 13 AND Y = 103 else
"100010011101" when X = 14 AND Y = 103 else
"100010011101" when X = 15 AND Y = 103 else
"100010011101" when X = 16 AND Y = 103 else
"100010011101" when X = 17 AND Y = 103 else
"100010011101" when X = 18 AND Y = 103 else
"100010011101" when X = 19 AND Y = 103 else
"110111011111" when X = 20 AND Y = 103 else
"110111011111" when X = 21 AND Y = 103 else
"110111011111" when X = 22 AND Y = 103 else
"110111011111" when X = 23 AND Y = 103 else
"110111011111" when X = 24 AND Y = 103 else
"110111011111" when X = 25 AND Y = 103 else
"110111011111" when X = 26 AND Y = 103 else
"110111011111" when X = 27 AND Y = 103 else
"110111011111" when X = 28 AND Y = 103 else
"110111011111" when X = 29 AND Y = 103 else
"110111011111" when X = 30 AND Y = 103 else
"110111011111" when X = 31 AND Y = 103 else
"110111011111" when X = 32 AND Y = 103 else
"110111011111" when X = 33 AND Y = 103 else
"110111011111" when X = 34 AND Y = 103 else
"110111011111" when X = 35 AND Y = 103 else
"110111011111" when X = 36 AND Y = 103 else
"110111011111" when X = 37 AND Y = 103 else
"110111011111" when X = 38 AND Y = 103 else
"110111011111" when X = 39 AND Y = 103 else
"110111011111" when X = 40 AND Y = 103 else
"110111011111" when X = 41 AND Y = 103 else
"110111011111" when X = 42 AND Y = 103 else
"110111011111" when X = 43 AND Y = 103 else
"110111011111" when X = 44 AND Y = 103 else
"110111011111" when X = 45 AND Y = 103 else
"110111011111" when X = 46 AND Y = 103 else
"110111011111" when X = 47 AND Y = 103 else
"110111011111" when X = 48 AND Y = 103 else
"110111011111" when X = 49 AND Y = 103 else
"110111011111" when X = 50 AND Y = 103 else
"110111011111" when X = 51 AND Y = 103 else
"110111011111" when X = 52 AND Y = 103 else
"110111011111" when X = 53 AND Y = 103 else
"110111011111" when X = 54 AND Y = 103 else
"110111011111" when X = 55 AND Y = 103 else
"110111011111" when X = 56 AND Y = 103 else
"110111011111" when X = 57 AND Y = 103 else
"110111011111" when X = 58 AND Y = 103 else
"110111011111" when X = 59 AND Y = 103 else
"110111011111" when X = 60 AND Y = 103 else
"110111011111" when X = 61 AND Y = 103 else
"110111011111" when X = 62 AND Y = 103 else
"110111011111" when X = 63 AND Y = 103 else
"110111011111" when X = 64 AND Y = 103 else
"110111011111" when X = 65 AND Y = 103 else
"110111011111" when X = 66 AND Y = 103 else
"110111011111" when X = 67 AND Y = 103 else
"110111011111" when X = 68 AND Y = 103 else
"110111011111" when X = 69 AND Y = 103 else
"111111111111" when X = 70 AND Y = 103 else
"111111111111" when X = 71 AND Y = 103 else
"111111111111" when X = 72 AND Y = 103 else
"111111111111" when X = 73 AND Y = 103 else
"111111111111" when X = 74 AND Y = 103 else
"111111111111" when X = 75 AND Y = 103 else
"111111111111" when X = 76 AND Y = 103 else
"111111111111" when X = 77 AND Y = 103 else
"111111111111" when X = 78 AND Y = 103 else
"111111111111" when X = 79 AND Y = 103 else
"111111111111" when X = 80 AND Y = 103 else
"111111111111" when X = 81 AND Y = 103 else
"111111111111" when X = 82 AND Y = 103 else
"111111111111" when X = 83 AND Y = 103 else
"111111111111" when X = 84 AND Y = 103 else
"111111111111" when X = 85 AND Y = 103 else
"111111111111" when X = 86 AND Y = 103 else
"111111111111" when X = 87 AND Y = 103 else
"111111111111" when X = 88 AND Y = 103 else
"111111111111" when X = 89 AND Y = 103 else
"111111111111" when X = 90 AND Y = 103 else
"111111111111" when X = 91 AND Y = 103 else
"111111111111" when X = 92 AND Y = 103 else
"111111111111" when X = 93 AND Y = 103 else
"111111111111" when X = 94 AND Y = 103 else
"111111111111" when X = 95 AND Y = 103 else
"111111111111" when X = 96 AND Y = 103 else
"111111111111" when X = 97 AND Y = 103 else
"111111111111" when X = 98 AND Y = 103 else
"111111111111" when X = 99 AND Y = 103 else
"111111111111" when X = 100 AND Y = 103 else
"111111111111" when X = 101 AND Y = 103 else
"111111111111" when X = 102 AND Y = 103 else
"111111111111" when X = 103 AND Y = 103 else
"111111111111" when X = 104 AND Y = 103 else
"111111111111" when X = 105 AND Y = 103 else
"111111111111" when X = 106 AND Y = 103 else
"111111111111" when X = 107 AND Y = 103 else
"111111111111" when X = 108 AND Y = 103 else
"111111111111" when X = 109 AND Y = 103 else
"111111111111" when X = 110 AND Y = 103 else
"111111111111" when X = 111 AND Y = 103 else
"111111111111" when X = 112 AND Y = 103 else
"111111111111" when X = 113 AND Y = 103 else
"111111111111" when X = 114 AND Y = 103 else
"111111111111" when X = 115 AND Y = 103 else
"111111111111" when X = 116 AND Y = 103 else
"111111111111" when X = 117 AND Y = 103 else
"111111111111" when X = 118 AND Y = 103 else
"111111111111" when X = 119 AND Y = 103 else
"111111111111" when X = 120 AND Y = 103 else
"111111111111" when X = 121 AND Y = 103 else
"111111111111" when X = 122 AND Y = 103 else
"111111111111" when X = 123 AND Y = 103 else
"111111111111" when X = 124 AND Y = 103 else
"111111111111" when X = 125 AND Y = 103 else
"111111111111" when X = 126 AND Y = 103 else
"111111111111" when X = 127 AND Y = 103 else
"111111111111" when X = 128 AND Y = 103 else
"111111111111" when X = 129 AND Y = 103 else
"111111111111" when X = 130 AND Y = 103 else
"111111111111" when X = 131 AND Y = 103 else
"111111111111" when X = 132 AND Y = 103 else
"111111111111" when X = 133 AND Y = 103 else
"111111111111" when X = 134 AND Y = 103 else
"111111111111" when X = 135 AND Y = 103 else
"111111111111" when X = 136 AND Y = 103 else
"111111111111" when X = 137 AND Y = 103 else
"111111111111" when X = 138 AND Y = 103 else
"111111111111" when X = 139 AND Y = 103 else
"111111111111" when X = 140 AND Y = 103 else
"111111111111" when X = 141 AND Y = 103 else
"111111111111" when X = 142 AND Y = 103 else
"111111111111" when X = 143 AND Y = 103 else
"111111111111" when X = 144 AND Y = 103 else
"111111111111" when X = 145 AND Y = 103 else
"111111111111" when X = 146 AND Y = 103 else
"111111111111" when X = 147 AND Y = 103 else
"111111111111" when X = 148 AND Y = 103 else
"111111111111" when X = 149 AND Y = 103 else
"111111111111" when X = 150 AND Y = 103 else
"111111111111" when X = 151 AND Y = 103 else
"111111111111" when X = 152 AND Y = 103 else
"111111111111" when X = 153 AND Y = 103 else
"111111111111" when X = 154 AND Y = 103 else
"111111111111" when X = 155 AND Y = 103 else
"111111111111" when X = 156 AND Y = 103 else
"111111111111" when X = 157 AND Y = 103 else
"111111111111" when X = 158 AND Y = 103 else
"111111111111" when X = 159 AND Y = 103 else
"110111011111" when X = 160 AND Y = 103 else
"110111011111" when X = 161 AND Y = 103 else
"110111011111" when X = 162 AND Y = 103 else
"110111011111" when X = 163 AND Y = 103 else
"110111011111" when X = 164 AND Y = 103 else
"110111011111" when X = 165 AND Y = 103 else
"110111011111" when X = 166 AND Y = 103 else
"110111011111" when X = 167 AND Y = 103 else
"110111011111" when X = 168 AND Y = 103 else
"110111011111" when X = 169 AND Y = 103 else
"110111011111" when X = 170 AND Y = 103 else
"110111011111" when X = 171 AND Y = 103 else
"110111011111" when X = 172 AND Y = 103 else
"110111011111" when X = 173 AND Y = 103 else
"110111011111" when X = 174 AND Y = 103 else
"110111011111" when X = 175 AND Y = 103 else
"110111011111" when X = 176 AND Y = 103 else
"110111011111" when X = 177 AND Y = 103 else
"110111011111" when X = 178 AND Y = 103 else
"110111011111" when X = 179 AND Y = 103 else
"110111011111" when X = 180 AND Y = 103 else
"110111011111" when X = 181 AND Y = 103 else
"110111011111" when X = 182 AND Y = 103 else
"110111011111" when X = 183 AND Y = 103 else
"110111011111" when X = 184 AND Y = 103 else
"110111011111" when X = 185 AND Y = 103 else
"110111011111" when X = 186 AND Y = 103 else
"110111011111" when X = 187 AND Y = 103 else
"110111011111" when X = 188 AND Y = 103 else
"110111011111" when X = 189 AND Y = 103 else
"110111011111" when X = 190 AND Y = 103 else
"110111011111" when X = 191 AND Y = 103 else
"110111011111" when X = 192 AND Y = 103 else
"110111011111" when X = 193 AND Y = 103 else
"110111011111" when X = 194 AND Y = 103 else
"110111011111" when X = 195 AND Y = 103 else
"110111011111" when X = 196 AND Y = 103 else
"110111011111" when X = 197 AND Y = 103 else
"110111011111" when X = 198 AND Y = 103 else
"110111011111" when X = 199 AND Y = 103 else
"110111011111" when X = 200 AND Y = 103 else
"110111011111" when X = 201 AND Y = 103 else
"110111011111" when X = 202 AND Y = 103 else
"110111011111" when X = 203 AND Y = 103 else
"110111011111" when X = 204 AND Y = 103 else
"110111011111" when X = 205 AND Y = 103 else
"110111011111" when X = 206 AND Y = 103 else
"110111011111" when X = 207 AND Y = 103 else
"110111011111" when X = 208 AND Y = 103 else
"110111011111" when X = 209 AND Y = 103 else
"110111011111" when X = 210 AND Y = 103 else
"110111011111" when X = 211 AND Y = 103 else
"110111011111" when X = 212 AND Y = 103 else
"110111011111" when X = 213 AND Y = 103 else
"110111011111" when X = 214 AND Y = 103 else
"111111111111" when X = 215 AND Y = 103 else
"111111111111" when X = 216 AND Y = 103 else
"111111111111" when X = 217 AND Y = 103 else
"111111111111" when X = 218 AND Y = 103 else
"111111111111" when X = 219 AND Y = 103 else
"111111111111" when X = 220 AND Y = 103 else
"111111111111" when X = 221 AND Y = 103 else
"111111111111" when X = 222 AND Y = 103 else
"111111111111" when X = 223 AND Y = 103 else
"111111111111" when X = 224 AND Y = 103 else
"111111111111" when X = 225 AND Y = 103 else
"111111111111" when X = 226 AND Y = 103 else
"111111111111" when X = 227 AND Y = 103 else
"111111111111" when X = 228 AND Y = 103 else
"111111111111" when X = 229 AND Y = 103 else
"111111111111" when X = 230 AND Y = 103 else
"111111111111" when X = 231 AND Y = 103 else
"111111111111" when X = 232 AND Y = 103 else
"111111111111" when X = 233 AND Y = 103 else
"111111111111" when X = 234 AND Y = 103 else
"111111111111" when X = 235 AND Y = 103 else
"111111111111" when X = 236 AND Y = 103 else
"111111111111" when X = 237 AND Y = 103 else
"111111111111" when X = 238 AND Y = 103 else
"111111111111" when X = 239 AND Y = 103 else
"110111011111" when X = 240 AND Y = 103 else
"110111011111" when X = 241 AND Y = 103 else
"110111011111" when X = 242 AND Y = 103 else
"110111011111" when X = 243 AND Y = 103 else
"110111011111" when X = 244 AND Y = 103 else
"110111011111" when X = 245 AND Y = 103 else
"110111011111" when X = 246 AND Y = 103 else
"110111011111" when X = 247 AND Y = 103 else
"110111011111" when X = 248 AND Y = 103 else
"110111011111" when X = 249 AND Y = 103 else
"111111111111" when X = 250 AND Y = 103 else
"111111111111" when X = 251 AND Y = 103 else
"111111111111" when X = 252 AND Y = 103 else
"111111111111" when X = 253 AND Y = 103 else
"111111111111" when X = 254 AND Y = 103 else
"111111111111" when X = 255 AND Y = 103 else
"111111111111" when X = 256 AND Y = 103 else
"111111111111" when X = 257 AND Y = 103 else
"111111111111" when X = 258 AND Y = 103 else
"111111111111" when X = 259 AND Y = 103 else
"111111111111" when X = 260 AND Y = 103 else
"111111111111" when X = 261 AND Y = 103 else
"111111111111" when X = 262 AND Y = 103 else
"111111111111" when X = 263 AND Y = 103 else
"111111111111" when X = 264 AND Y = 103 else
"111111111111" when X = 265 AND Y = 103 else
"111111111111" when X = 266 AND Y = 103 else
"111111111111" when X = 267 AND Y = 103 else
"111111111111" when X = 268 AND Y = 103 else
"111111111111" when X = 269 AND Y = 103 else
"111111111111" when X = 270 AND Y = 103 else
"111111111111" when X = 271 AND Y = 103 else
"111111111111" when X = 272 AND Y = 103 else
"111111111111" when X = 273 AND Y = 103 else
"111111111111" when X = 274 AND Y = 103 else
"110111011111" when X = 275 AND Y = 103 else
"110111011111" when X = 276 AND Y = 103 else
"110111011111" when X = 277 AND Y = 103 else
"110111011111" when X = 278 AND Y = 103 else
"110111011111" when X = 279 AND Y = 103 else
"111111111111" when X = 280 AND Y = 103 else
"111111111111" when X = 281 AND Y = 103 else
"111111111111" when X = 282 AND Y = 103 else
"111111111111" when X = 283 AND Y = 103 else
"111111111111" when X = 284 AND Y = 103 else
"111111111111" when X = 285 AND Y = 103 else
"111111111111" when X = 286 AND Y = 103 else
"111111111111" when X = 287 AND Y = 103 else
"111111111111" when X = 288 AND Y = 103 else
"111111111111" when X = 289 AND Y = 103 else
"111111111111" when X = 290 AND Y = 103 else
"111111111111" when X = 291 AND Y = 103 else
"111111111111" when X = 292 AND Y = 103 else
"111111111111" when X = 293 AND Y = 103 else
"111111111111" when X = 294 AND Y = 103 else
"111111111111" when X = 295 AND Y = 103 else
"111111111111" when X = 296 AND Y = 103 else
"111111111111" when X = 297 AND Y = 103 else
"111111111111" when X = 298 AND Y = 103 else
"111111111111" when X = 299 AND Y = 103 else
"111111111111" when X = 300 AND Y = 103 else
"111111111111" when X = 301 AND Y = 103 else
"111111111111" when X = 302 AND Y = 103 else
"111111111111" when X = 303 AND Y = 103 else
"111111111111" when X = 304 AND Y = 103 else
"110111011111" when X = 305 AND Y = 103 else
"110111011111" when X = 306 AND Y = 103 else
"110111011111" when X = 307 AND Y = 103 else
"110111011111" when X = 308 AND Y = 103 else
"110111011111" when X = 309 AND Y = 103 else
"110111011111" when X = 310 AND Y = 103 else
"110111011111" when X = 311 AND Y = 103 else
"110111011111" when X = 312 AND Y = 103 else
"110111011111" when X = 313 AND Y = 103 else
"110111011111" when X = 314 AND Y = 103 else
"110111011111" when X = 315 AND Y = 103 else
"110111011111" when X = 316 AND Y = 103 else
"110111011111" when X = 317 AND Y = 103 else
"110111011111" when X = 318 AND Y = 103 else
"110111011111" when X = 319 AND Y = 103 else
"110111011111" when X = 320 AND Y = 103 else
"110111011111" when X = 321 AND Y = 103 else
"110111011111" when X = 322 AND Y = 103 else
"110111011111" when X = 323 AND Y = 103 else
"110111011111" when X = 324 AND Y = 103 else
"100010011101" when X = 0 AND Y = 104 else
"100010011101" when X = 1 AND Y = 104 else
"100010011101" when X = 2 AND Y = 104 else
"100010011101" when X = 3 AND Y = 104 else
"100010011101" when X = 4 AND Y = 104 else
"100010011101" when X = 5 AND Y = 104 else
"100010011101" when X = 6 AND Y = 104 else
"100010011101" when X = 7 AND Y = 104 else
"100010011101" when X = 8 AND Y = 104 else
"100010011101" when X = 9 AND Y = 104 else
"100010011101" when X = 10 AND Y = 104 else
"100010011101" when X = 11 AND Y = 104 else
"100010011101" when X = 12 AND Y = 104 else
"100010011101" when X = 13 AND Y = 104 else
"100010011101" when X = 14 AND Y = 104 else
"100010011101" when X = 15 AND Y = 104 else
"100010011101" when X = 16 AND Y = 104 else
"100010011101" when X = 17 AND Y = 104 else
"100010011101" when X = 18 AND Y = 104 else
"100010011101" when X = 19 AND Y = 104 else
"110111011111" when X = 20 AND Y = 104 else
"110111011111" when X = 21 AND Y = 104 else
"110111011111" when X = 22 AND Y = 104 else
"110111011111" when X = 23 AND Y = 104 else
"110111011111" when X = 24 AND Y = 104 else
"110111011111" when X = 25 AND Y = 104 else
"110111011111" when X = 26 AND Y = 104 else
"110111011111" when X = 27 AND Y = 104 else
"110111011111" when X = 28 AND Y = 104 else
"110111011111" when X = 29 AND Y = 104 else
"110111011111" when X = 30 AND Y = 104 else
"110111011111" when X = 31 AND Y = 104 else
"110111011111" when X = 32 AND Y = 104 else
"110111011111" when X = 33 AND Y = 104 else
"110111011111" when X = 34 AND Y = 104 else
"110111011111" when X = 35 AND Y = 104 else
"110111011111" when X = 36 AND Y = 104 else
"110111011111" when X = 37 AND Y = 104 else
"110111011111" when X = 38 AND Y = 104 else
"110111011111" when X = 39 AND Y = 104 else
"110111011111" when X = 40 AND Y = 104 else
"110111011111" when X = 41 AND Y = 104 else
"110111011111" when X = 42 AND Y = 104 else
"110111011111" when X = 43 AND Y = 104 else
"110111011111" when X = 44 AND Y = 104 else
"110111011111" when X = 45 AND Y = 104 else
"110111011111" when X = 46 AND Y = 104 else
"110111011111" when X = 47 AND Y = 104 else
"110111011111" when X = 48 AND Y = 104 else
"110111011111" when X = 49 AND Y = 104 else
"110111011111" when X = 50 AND Y = 104 else
"110111011111" when X = 51 AND Y = 104 else
"110111011111" when X = 52 AND Y = 104 else
"110111011111" when X = 53 AND Y = 104 else
"110111011111" when X = 54 AND Y = 104 else
"110111011111" when X = 55 AND Y = 104 else
"110111011111" when X = 56 AND Y = 104 else
"110111011111" when X = 57 AND Y = 104 else
"110111011111" when X = 58 AND Y = 104 else
"110111011111" when X = 59 AND Y = 104 else
"110111011111" when X = 60 AND Y = 104 else
"110111011111" when X = 61 AND Y = 104 else
"110111011111" when X = 62 AND Y = 104 else
"110111011111" when X = 63 AND Y = 104 else
"110111011111" when X = 64 AND Y = 104 else
"110111011111" when X = 65 AND Y = 104 else
"110111011111" when X = 66 AND Y = 104 else
"110111011111" when X = 67 AND Y = 104 else
"110111011111" when X = 68 AND Y = 104 else
"110111011111" when X = 69 AND Y = 104 else
"111111111111" when X = 70 AND Y = 104 else
"111111111111" when X = 71 AND Y = 104 else
"111111111111" when X = 72 AND Y = 104 else
"111111111111" when X = 73 AND Y = 104 else
"111111111111" when X = 74 AND Y = 104 else
"111111111111" when X = 75 AND Y = 104 else
"111111111111" when X = 76 AND Y = 104 else
"111111111111" when X = 77 AND Y = 104 else
"111111111111" when X = 78 AND Y = 104 else
"111111111111" when X = 79 AND Y = 104 else
"111111111111" when X = 80 AND Y = 104 else
"111111111111" when X = 81 AND Y = 104 else
"111111111111" when X = 82 AND Y = 104 else
"111111111111" when X = 83 AND Y = 104 else
"111111111111" when X = 84 AND Y = 104 else
"111111111111" when X = 85 AND Y = 104 else
"111111111111" when X = 86 AND Y = 104 else
"111111111111" when X = 87 AND Y = 104 else
"111111111111" when X = 88 AND Y = 104 else
"111111111111" when X = 89 AND Y = 104 else
"111111111111" when X = 90 AND Y = 104 else
"111111111111" when X = 91 AND Y = 104 else
"111111111111" when X = 92 AND Y = 104 else
"111111111111" when X = 93 AND Y = 104 else
"111111111111" when X = 94 AND Y = 104 else
"111111111111" when X = 95 AND Y = 104 else
"111111111111" when X = 96 AND Y = 104 else
"111111111111" when X = 97 AND Y = 104 else
"111111111111" when X = 98 AND Y = 104 else
"111111111111" when X = 99 AND Y = 104 else
"111111111111" when X = 100 AND Y = 104 else
"111111111111" when X = 101 AND Y = 104 else
"111111111111" when X = 102 AND Y = 104 else
"111111111111" when X = 103 AND Y = 104 else
"111111111111" when X = 104 AND Y = 104 else
"111111111111" when X = 105 AND Y = 104 else
"111111111111" when X = 106 AND Y = 104 else
"111111111111" when X = 107 AND Y = 104 else
"111111111111" when X = 108 AND Y = 104 else
"111111111111" when X = 109 AND Y = 104 else
"111111111111" when X = 110 AND Y = 104 else
"111111111111" when X = 111 AND Y = 104 else
"111111111111" when X = 112 AND Y = 104 else
"111111111111" when X = 113 AND Y = 104 else
"111111111111" when X = 114 AND Y = 104 else
"111111111111" when X = 115 AND Y = 104 else
"111111111111" when X = 116 AND Y = 104 else
"111111111111" when X = 117 AND Y = 104 else
"111111111111" when X = 118 AND Y = 104 else
"111111111111" when X = 119 AND Y = 104 else
"111111111111" when X = 120 AND Y = 104 else
"111111111111" when X = 121 AND Y = 104 else
"111111111111" when X = 122 AND Y = 104 else
"111111111111" when X = 123 AND Y = 104 else
"111111111111" when X = 124 AND Y = 104 else
"111111111111" when X = 125 AND Y = 104 else
"111111111111" when X = 126 AND Y = 104 else
"111111111111" when X = 127 AND Y = 104 else
"111111111111" when X = 128 AND Y = 104 else
"111111111111" when X = 129 AND Y = 104 else
"111111111111" when X = 130 AND Y = 104 else
"111111111111" when X = 131 AND Y = 104 else
"111111111111" when X = 132 AND Y = 104 else
"111111111111" when X = 133 AND Y = 104 else
"111111111111" when X = 134 AND Y = 104 else
"111111111111" when X = 135 AND Y = 104 else
"111111111111" when X = 136 AND Y = 104 else
"111111111111" when X = 137 AND Y = 104 else
"111111111111" when X = 138 AND Y = 104 else
"111111111111" when X = 139 AND Y = 104 else
"111111111111" when X = 140 AND Y = 104 else
"111111111111" when X = 141 AND Y = 104 else
"111111111111" when X = 142 AND Y = 104 else
"111111111111" when X = 143 AND Y = 104 else
"111111111111" when X = 144 AND Y = 104 else
"111111111111" when X = 145 AND Y = 104 else
"111111111111" when X = 146 AND Y = 104 else
"111111111111" when X = 147 AND Y = 104 else
"111111111111" when X = 148 AND Y = 104 else
"111111111111" when X = 149 AND Y = 104 else
"111111111111" when X = 150 AND Y = 104 else
"111111111111" when X = 151 AND Y = 104 else
"111111111111" when X = 152 AND Y = 104 else
"111111111111" when X = 153 AND Y = 104 else
"111111111111" when X = 154 AND Y = 104 else
"111111111111" when X = 155 AND Y = 104 else
"111111111111" when X = 156 AND Y = 104 else
"111111111111" when X = 157 AND Y = 104 else
"111111111111" when X = 158 AND Y = 104 else
"111111111111" when X = 159 AND Y = 104 else
"110111011111" when X = 160 AND Y = 104 else
"110111011111" when X = 161 AND Y = 104 else
"110111011111" when X = 162 AND Y = 104 else
"110111011111" when X = 163 AND Y = 104 else
"110111011111" when X = 164 AND Y = 104 else
"110111011111" when X = 165 AND Y = 104 else
"110111011111" when X = 166 AND Y = 104 else
"110111011111" when X = 167 AND Y = 104 else
"110111011111" when X = 168 AND Y = 104 else
"110111011111" when X = 169 AND Y = 104 else
"110111011111" when X = 170 AND Y = 104 else
"110111011111" when X = 171 AND Y = 104 else
"110111011111" when X = 172 AND Y = 104 else
"110111011111" when X = 173 AND Y = 104 else
"110111011111" when X = 174 AND Y = 104 else
"110111011111" when X = 175 AND Y = 104 else
"110111011111" when X = 176 AND Y = 104 else
"110111011111" when X = 177 AND Y = 104 else
"110111011111" when X = 178 AND Y = 104 else
"110111011111" when X = 179 AND Y = 104 else
"110111011111" when X = 180 AND Y = 104 else
"110111011111" when X = 181 AND Y = 104 else
"110111011111" when X = 182 AND Y = 104 else
"110111011111" when X = 183 AND Y = 104 else
"110111011111" when X = 184 AND Y = 104 else
"110111011111" when X = 185 AND Y = 104 else
"110111011111" when X = 186 AND Y = 104 else
"110111011111" when X = 187 AND Y = 104 else
"110111011111" when X = 188 AND Y = 104 else
"110111011111" when X = 189 AND Y = 104 else
"110111011111" when X = 190 AND Y = 104 else
"110111011111" when X = 191 AND Y = 104 else
"110111011111" when X = 192 AND Y = 104 else
"110111011111" when X = 193 AND Y = 104 else
"110111011111" when X = 194 AND Y = 104 else
"110111011111" when X = 195 AND Y = 104 else
"110111011111" when X = 196 AND Y = 104 else
"110111011111" when X = 197 AND Y = 104 else
"110111011111" when X = 198 AND Y = 104 else
"110111011111" when X = 199 AND Y = 104 else
"110111011111" when X = 200 AND Y = 104 else
"110111011111" when X = 201 AND Y = 104 else
"110111011111" when X = 202 AND Y = 104 else
"110111011111" when X = 203 AND Y = 104 else
"110111011111" when X = 204 AND Y = 104 else
"110111011111" when X = 205 AND Y = 104 else
"110111011111" when X = 206 AND Y = 104 else
"110111011111" when X = 207 AND Y = 104 else
"110111011111" when X = 208 AND Y = 104 else
"110111011111" when X = 209 AND Y = 104 else
"110111011111" when X = 210 AND Y = 104 else
"110111011111" when X = 211 AND Y = 104 else
"110111011111" when X = 212 AND Y = 104 else
"110111011111" when X = 213 AND Y = 104 else
"110111011111" when X = 214 AND Y = 104 else
"111111111111" when X = 215 AND Y = 104 else
"111111111111" when X = 216 AND Y = 104 else
"111111111111" when X = 217 AND Y = 104 else
"111111111111" when X = 218 AND Y = 104 else
"111111111111" when X = 219 AND Y = 104 else
"111111111111" when X = 220 AND Y = 104 else
"111111111111" when X = 221 AND Y = 104 else
"111111111111" when X = 222 AND Y = 104 else
"111111111111" when X = 223 AND Y = 104 else
"111111111111" when X = 224 AND Y = 104 else
"111111111111" when X = 225 AND Y = 104 else
"111111111111" when X = 226 AND Y = 104 else
"111111111111" when X = 227 AND Y = 104 else
"111111111111" when X = 228 AND Y = 104 else
"111111111111" when X = 229 AND Y = 104 else
"111111111111" when X = 230 AND Y = 104 else
"111111111111" when X = 231 AND Y = 104 else
"111111111111" when X = 232 AND Y = 104 else
"111111111111" when X = 233 AND Y = 104 else
"111111111111" when X = 234 AND Y = 104 else
"111111111111" when X = 235 AND Y = 104 else
"111111111111" when X = 236 AND Y = 104 else
"111111111111" when X = 237 AND Y = 104 else
"111111111111" when X = 238 AND Y = 104 else
"111111111111" when X = 239 AND Y = 104 else
"110111011111" when X = 240 AND Y = 104 else
"110111011111" when X = 241 AND Y = 104 else
"110111011111" when X = 242 AND Y = 104 else
"110111011111" when X = 243 AND Y = 104 else
"110111011111" when X = 244 AND Y = 104 else
"110111011111" when X = 245 AND Y = 104 else
"110111011111" when X = 246 AND Y = 104 else
"110111011111" when X = 247 AND Y = 104 else
"110111011111" when X = 248 AND Y = 104 else
"110111011111" when X = 249 AND Y = 104 else
"111111111111" when X = 250 AND Y = 104 else
"111111111111" when X = 251 AND Y = 104 else
"111111111111" when X = 252 AND Y = 104 else
"111111111111" when X = 253 AND Y = 104 else
"111111111111" when X = 254 AND Y = 104 else
"111111111111" when X = 255 AND Y = 104 else
"111111111111" when X = 256 AND Y = 104 else
"111111111111" when X = 257 AND Y = 104 else
"111111111111" when X = 258 AND Y = 104 else
"111111111111" when X = 259 AND Y = 104 else
"111111111111" when X = 260 AND Y = 104 else
"111111111111" when X = 261 AND Y = 104 else
"111111111111" when X = 262 AND Y = 104 else
"111111111111" when X = 263 AND Y = 104 else
"111111111111" when X = 264 AND Y = 104 else
"111111111111" when X = 265 AND Y = 104 else
"111111111111" when X = 266 AND Y = 104 else
"111111111111" when X = 267 AND Y = 104 else
"111111111111" when X = 268 AND Y = 104 else
"111111111111" when X = 269 AND Y = 104 else
"111111111111" when X = 270 AND Y = 104 else
"111111111111" when X = 271 AND Y = 104 else
"111111111111" when X = 272 AND Y = 104 else
"111111111111" when X = 273 AND Y = 104 else
"111111111111" when X = 274 AND Y = 104 else
"110111011111" when X = 275 AND Y = 104 else
"110111011111" when X = 276 AND Y = 104 else
"110111011111" when X = 277 AND Y = 104 else
"110111011111" when X = 278 AND Y = 104 else
"110111011111" when X = 279 AND Y = 104 else
"111111111111" when X = 280 AND Y = 104 else
"111111111111" when X = 281 AND Y = 104 else
"111111111111" when X = 282 AND Y = 104 else
"111111111111" when X = 283 AND Y = 104 else
"111111111111" when X = 284 AND Y = 104 else
"111111111111" when X = 285 AND Y = 104 else
"111111111111" when X = 286 AND Y = 104 else
"111111111111" when X = 287 AND Y = 104 else
"111111111111" when X = 288 AND Y = 104 else
"111111111111" when X = 289 AND Y = 104 else
"111111111111" when X = 290 AND Y = 104 else
"111111111111" when X = 291 AND Y = 104 else
"111111111111" when X = 292 AND Y = 104 else
"111111111111" when X = 293 AND Y = 104 else
"111111111111" when X = 294 AND Y = 104 else
"111111111111" when X = 295 AND Y = 104 else
"111111111111" when X = 296 AND Y = 104 else
"111111111111" when X = 297 AND Y = 104 else
"111111111111" when X = 298 AND Y = 104 else
"111111111111" when X = 299 AND Y = 104 else
"111111111111" when X = 300 AND Y = 104 else
"111111111111" when X = 301 AND Y = 104 else
"111111111111" when X = 302 AND Y = 104 else
"111111111111" when X = 303 AND Y = 104 else
"111111111111" when X = 304 AND Y = 104 else
"110111011111" when X = 305 AND Y = 104 else
"110111011111" when X = 306 AND Y = 104 else
"110111011111" when X = 307 AND Y = 104 else
"110111011111" when X = 308 AND Y = 104 else
"110111011111" when X = 309 AND Y = 104 else
"110111011111" when X = 310 AND Y = 104 else
"110111011111" when X = 311 AND Y = 104 else
"110111011111" when X = 312 AND Y = 104 else
"110111011111" when X = 313 AND Y = 104 else
"110111011111" when X = 314 AND Y = 104 else
"110111011111" when X = 315 AND Y = 104 else
"110111011111" when X = 316 AND Y = 104 else
"110111011111" when X = 317 AND Y = 104 else
"110111011111" when X = 318 AND Y = 104 else
"110111011111" when X = 319 AND Y = 104 else
"110111011111" when X = 320 AND Y = 104 else
"110111011111" when X = 321 AND Y = 104 else
"110111011111" when X = 322 AND Y = 104 else
"110111011111" when X = 323 AND Y = 104 else
"110111011111" when X = 324 AND Y = 104 else
"100010011101" when X = 0 AND Y = 105 else
"100010011101" when X = 1 AND Y = 105 else
"100010011101" when X = 2 AND Y = 105 else
"100010011101" when X = 3 AND Y = 105 else
"100010011101" when X = 4 AND Y = 105 else
"100010011101" when X = 5 AND Y = 105 else
"100010011101" when X = 6 AND Y = 105 else
"100010011101" when X = 7 AND Y = 105 else
"100010011101" when X = 8 AND Y = 105 else
"100010011101" when X = 9 AND Y = 105 else
"100010011101" when X = 10 AND Y = 105 else
"100010011101" when X = 11 AND Y = 105 else
"100010011101" when X = 12 AND Y = 105 else
"100010011101" when X = 13 AND Y = 105 else
"100010011101" when X = 14 AND Y = 105 else
"100010011101" when X = 15 AND Y = 105 else
"100010011101" when X = 16 AND Y = 105 else
"100010011101" when X = 17 AND Y = 105 else
"100010011101" when X = 18 AND Y = 105 else
"100010011101" when X = 19 AND Y = 105 else
"100010011101" when X = 20 AND Y = 105 else
"100010011101" when X = 21 AND Y = 105 else
"100010011101" when X = 22 AND Y = 105 else
"100010011101" when X = 23 AND Y = 105 else
"100010011101" when X = 24 AND Y = 105 else
"110111011111" when X = 25 AND Y = 105 else
"110111011111" when X = 26 AND Y = 105 else
"110111011111" when X = 27 AND Y = 105 else
"110111011111" when X = 28 AND Y = 105 else
"110111011111" when X = 29 AND Y = 105 else
"110111011111" when X = 30 AND Y = 105 else
"110111011111" when X = 31 AND Y = 105 else
"110111011111" when X = 32 AND Y = 105 else
"110111011111" when X = 33 AND Y = 105 else
"110111011111" when X = 34 AND Y = 105 else
"110111011111" when X = 35 AND Y = 105 else
"110111011111" when X = 36 AND Y = 105 else
"110111011111" when X = 37 AND Y = 105 else
"110111011111" when X = 38 AND Y = 105 else
"110111011111" when X = 39 AND Y = 105 else
"110111011111" when X = 40 AND Y = 105 else
"110111011111" when X = 41 AND Y = 105 else
"110111011111" when X = 42 AND Y = 105 else
"110111011111" when X = 43 AND Y = 105 else
"110111011111" when X = 44 AND Y = 105 else
"110111011111" when X = 45 AND Y = 105 else
"110111011111" when X = 46 AND Y = 105 else
"110111011111" when X = 47 AND Y = 105 else
"110111011111" when X = 48 AND Y = 105 else
"110111011111" when X = 49 AND Y = 105 else
"110111011111" when X = 50 AND Y = 105 else
"110111011111" when X = 51 AND Y = 105 else
"110111011111" when X = 52 AND Y = 105 else
"110111011111" when X = 53 AND Y = 105 else
"110111011111" when X = 54 AND Y = 105 else
"110111011111" when X = 55 AND Y = 105 else
"110111011111" when X = 56 AND Y = 105 else
"110111011111" when X = 57 AND Y = 105 else
"110111011111" when X = 58 AND Y = 105 else
"110111011111" when X = 59 AND Y = 105 else
"110111011111" when X = 60 AND Y = 105 else
"110111011111" when X = 61 AND Y = 105 else
"110111011111" when X = 62 AND Y = 105 else
"110111011111" when X = 63 AND Y = 105 else
"110111011111" when X = 64 AND Y = 105 else
"110111011111" when X = 65 AND Y = 105 else
"110111011111" when X = 66 AND Y = 105 else
"110111011111" when X = 67 AND Y = 105 else
"110111011111" when X = 68 AND Y = 105 else
"110111011111" when X = 69 AND Y = 105 else
"111111111111" when X = 70 AND Y = 105 else
"111111111111" when X = 71 AND Y = 105 else
"111111111111" when X = 72 AND Y = 105 else
"111111111111" when X = 73 AND Y = 105 else
"111111111111" when X = 74 AND Y = 105 else
"111111111111" when X = 75 AND Y = 105 else
"111111111111" when X = 76 AND Y = 105 else
"111111111111" when X = 77 AND Y = 105 else
"111111111111" when X = 78 AND Y = 105 else
"111111111111" when X = 79 AND Y = 105 else
"111111111111" when X = 80 AND Y = 105 else
"111111111111" when X = 81 AND Y = 105 else
"111111111111" when X = 82 AND Y = 105 else
"111111111111" when X = 83 AND Y = 105 else
"111111111111" when X = 84 AND Y = 105 else
"111111111111" when X = 85 AND Y = 105 else
"111111111111" when X = 86 AND Y = 105 else
"111111111111" when X = 87 AND Y = 105 else
"111111111111" when X = 88 AND Y = 105 else
"111111111111" when X = 89 AND Y = 105 else
"111111111111" when X = 90 AND Y = 105 else
"111111111111" when X = 91 AND Y = 105 else
"111111111111" when X = 92 AND Y = 105 else
"111111111111" when X = 93 AND Y = 105 else
"111111111111" when X = 94 AND Y = 105 else
"111111111111" when X = 95 AND Y = 105 else
"111111111111" when X = 96 AND Y = 105 else
"111111111111" when X = 97 AND Y = 105 else
"111111111111" when X = 98 AND Y = 105 else
"111111111111" when X = 99 AND Y = 105 else
"111111111111" when X = 100 AND Y = 105 else
"111111111111" when X = 101 AND Y = 105 else
"111111111111" when X = 102 AND Y = 105 else
"111111111111" when X = 103 AND Y = 105 else
"111111111111" when X = 104 AND Y = 105 else
"111111111111" when X = 105 AND Y = 105 else
"111111111111" when X = 106 AND Y = 105 else
"111111111111" when X = 107 AND Y = 105 else
"111111111111" when X = 108 AND Y = 105 else
"111111111111" when X = 109 AND Y = 105 else
"111111111111" when X = 110 AND Y = 105 else
"111111111111" when X = 111 AND Y = 105 else
"111111111111" when X = 112 AND Y = 105 else
"111111111111" when X = 113 AND Y = 105 else
"111111111111" when X = 114 AND Y = 105 else
"111111111111" when X = 115 AND Y = 105 else
"111111111111" when X = 116 AND Y = 105 else
"111111111111" when X = 117 AND Y = 105 else
"111111111111" when X = 118 AND Y = 105 else
"111111111111" when X = 119 AND Y = 105 else
"111111111111" when X = 120 AND Y = 105 else
"111111111111" when X = 121 AND Y = 105 else
"111111111111" when X = 122 AND Y = 105 else
"111111111111" when X = 123 AND Y = 105 else
"111111111111" when X = 124 AND Y = 105 else
"111111111111" when X = 125 AND Y = 105 else
"111111111111" when X = 126 AND Y = 105 else
"111111111111" when X = 127 AND Y = 105 else
"111111111111" when X = 128 AND Y = 105 else
"111111111111" when X = 129 AND Y = 105 else
"111111111111" when X = 130 AND Y = 105 else
"111111111111" when X = 131 AND Y = 105 else
"111111111111" when X = 132 AND Y = 105 else
"111111111111" when X = 133 AND Y = 105 else
"111111111111" when X = 134 AND Y = 105 else
"111111111111" when X = 135 AND Y = 105 else
"111111111111" when X = 136 AND Y = 105 else
"111111111111" when X = 137 AND Y = 105 else
"111111111111" when X = 138 AND Y = 105 else
"111111111111" when X = 139 AND Y = 105 else
"111111111111" when X = 140 AND Y = 105 else
"111111111111" when X = 141 AND Y = 105 else
"111111111111" when X = 142 AND Y = 105 else
"111111111111" when X = 143 AND Y = 105 else
"111111111111" when X = 144 AND Y = 105 else
"111111111111" when X = 145 AND Y = 105 else
"111111111111" when X = 146 AND Y = 105 else
"111111111111" when X = 147 AND Y = 105 else
"111111111111" when X = 148 AND Y = 105 else
"111111111111" when X = 149 AND Y = 105 else
"111111111111" when X = 150 AND Y = 105 else
"111111111111" when X = 151 AND Y = 105 else
"111111111111" when X = 152 AND Y = 105 else
"111111111111" when X = 153 AND Y = 105 else
"111111111111" when X = 154 AND Y = 105 else
"111111111111" when X = 155 AND Y = 105 else
"111111111111" when X = 156 AND Y = 105 else
"111111111111" when X = 157 AND Y = 105 else
"111111111111" when X = 158 AND Y = 105 else
"111111111111" when X = 159 AND Y = 105 else
"110111011111" when X = 160 AND Y = 105 else
"110111011111" when X = 161 AND Y = 105 else
"110111011111" when X = 162 AND Y = 105 else
"110111011111" when X = 163 AND Y = 105 else
"110111011111" when X = 164 AND Y = 105 else
"110111011111" when X = 165 AND Y = 105 else
"110111011111" when X = 166 AND Y = 105 else
"110111011111" when X = 167 AND Y = 105 else
"110111011111" when X = 168 AND Y = 105 else
"110111011111" when X = 169 AND Y = 105 else
"110111011111" when X = 170 AND Y = 105 else
"110111011111" when X = 171 AND Y = 105 else
"110111011111" when X = 172 AND Y = 105 else
"110111011111" when X = 173 AND Y = 105 else
"110111011111" when X = 174 AND Y = 105 else
"110111011111" when X = 175 AND Y = 105 else
"110111011111" when X = 176 AND Y = 105 else
"110111011111" when X = 177 AND Y = 105 else
"110111011111" when X = 178 AND Y = 105 else
"110111011111" when X = 179 AND Y = 105 else
"110111011111" when X = 180 AND Y = 105 else
"110111011111" when X = 181 AND Y = 105 else
"110111011111" when X = 182 AND Y = 105 else
"110111011111" when X = 183 AND Y = 105 else
"110111011111" when X = 184 AND Y = 105 else
"110111011111" when X = 185 AND Y = 105 else
"110111011111" when X = 186 AND Y = 105 else
"110111011111" when X = 187 AND Y = 105 else
"110111011111" when X = 188 AND Y = 105 else
"110111011111" when X = 189 AND Y = 105 else
"110111011111" when X = 190 AND Y = 105 else
"110111011111" when X = 191 AND Y = 105 else
"110111011111" when X = 192 AND Y = 105 else
"110111011111" when X = 193 AND Y = 105 else
"110111011111" when X = 194 AND Y = 105 else
"110111011111" when X = 195 AND Y = 105 else
"110111011111" when X = 196 AND Y = 105 else
"110111011111" when X = 197 AND Y = 105 else
"110111011111" when X = 198 AND Y = 105 else
"110111011111" when X = 199 AND Y = 105 else
"110111011111" when X = 200 AND Y = 105 else
"110111011111" when X = 201 AND Y = 105 else
"110111011111" when X = 202 AND Y = 105 else
"110111011111" when X = 203 AND Y = 105 else
"110111011111" when X = 204 AND Y = 105 else
"111111111111" when X = 205 AND Y = 105 else
"111111111111" when X = 206 AND Y = 105 else
"111111111111" when X = 207 AND Y = 105 else
"111111111111" when X = 208 AND Y = 105 else
"111111111111" when X = 209 AND Y = 105 else
"111111111111" when X = 210 AND Y = 105 else
"111111111111" when X = 211 AND Y = 105 else
"111111111111" when X = 212 AND Y = 105 else
"111111111111" when X = 213 AND Y = 105 else
"111111111111" when X = 214 AND Y = 105 else
"110111011111" when X = 215 AND Y = 105 else
"110111011111" when X = 216 AND Y = 105 else
"110111011111" when X = 217 AND Y = 105 else
"110111011111" when X = 218 AND Y = 105 else
"110111011111" when X = 219 AND Y = 105 else
"110111011111" when X = 220 AND Y = 105 else
"110111011111" when X = 221 AND Y = 105 else
"110111011111" when X = 222 AND Y = 105 else
"110111011111" when X = 223 AND Y = 105 else
"110111011111" when X = 224 AND Y = 105 else
"110111011111" when X = 225 AND Y = 105 else
"110111011111" when X = 226 AND Y = 105 else
"110111011111" when X = 227 AND Y = 105 else
"110111011111" when X = 228 AND Y = 105 else
"110111011111" when X = 229 AND Y = 105 else
"110111011111" when X = 230 AND Y = 105 else
"110111011111" when X = 231 AND Y = 105 else
"110111011111" when X = 232 AND Y = 105 else
"110111011111" when X = 233 AND Y = 105 else
"110111011111" when X = 234 AND Y = 105 else
"110111011111" when X = 235 AND Y = 105 else
"110111011111" when X = 236 AND Y = 105 else
"110111011111" when X = 237 AND Y = 105 else
"110111011111" when X = 238 AND Y = 105 else
"110111011111" when X = 239 AND Y = 105 else
"110111011111" when X = 240 AND Y = 105 else
"110111011111" when X = 241 AND Y = 105 else
"110111011111" when X = 242 AND Y = 105 else
"110111011111" when X = 243 AND Y = 105 else
"110111011111" when X = 244 AND Y = 105 else
"110111011111" when X = 245 AND Y = 105 else
"110111011111" when X = 246 AND Y = 105 else
"110111011111" when X = 247 AND Y = 105 else
"110111011111" when X = 248 AND Y = 105 else
"110111011111" when X = 249 AND Y = 105 else
"110111011111" when X = 250 AND Y = 105 else
"110111011111" when X = 251 AND Y = 105 else
"110111011111" when X = 252 AND Y = 105 else
"110111011111" when X = 253 AND Y = 105 else
"110111011111" when X = 254 AND Y = 105 else
"110111011111" when X = 255 AND Y = 105 else
"110111011111" when X = 256 AND Y = 105 else
"110111011111" when X = 257 AND Y = 105 else
"110111011111" when X = 258 AND Y = 105 else
"110111011111" when X = 259 AND Y = 105 else
"110111011111" when X = 260 AND Y = 105 else
"110111011111" when X = 261 AND Y = 105 else
"110111011111" when X = 262 AND Y = 105 else
"110111011111" when X = 263 AND Y = 105 else
"110111011111" when X = 264 AND Y = 105 else
"110111011111" when X = 265 AND Y = 105 else
"110111011111" when X = 266 AND Y = 105 else
"110111011111" when X = 267 AND Y = 105 else
"110111011111" when X = 268 AND Y = 105 else
"110111011111" when X = 269 AND Y = 105 else
"110111011111" when X = 270 AND Y = 105 else
"110111011111" when X = 271 AND Y = 105 else
"110111011111" when X = 272 AND Y = 105 else
"110111011111" when X = 273 AND Y = 105 else
"110111011111" when X = 274 AND Y = 105 else
"110111011111" when X = 275 AND Y = 105 else
"110111011111" when X = 276 AND Y = 105 else
"110111011111" when X = 277 AND Y = 105 else
"110111011111" when X = 278 AND Y = 105 else
"110111011111" when X = 279 AND Y = 105 else
"111111111111" when X = 280 AND Y = 105 else
"111111111111" when X = 281 AND Y = 105 else
"111111111111" when X = 282 AND Y = 105 else
"111111111111" when X = 283 AND Y = 105 else
"111111111111" when X = 284 AND Y = 105 else
"111111111111" when X = 285 AND Y = 105 else
"111111111111" when X = 286 AND Y = 105 else
"111111111111" when X = 287 AND Y = 105 else
"111111111111" when X = 288 AND Y = 105 else
"111111111111" when X = 289 AND Y = 105 else
"111111111111" when X = 290 AND Y = 105 else
"111111111111" when X = 291 AND Y = 105 else
"111111111111" when X = 292 AND Y = 105 else
"111111111111" when X = 293 AND Y = 105 else
"111111111111" when X = 294 AND Y = 105 else
"111111111111" when X = 295 AND Y = 105 else
"111111111111" when X = 296 AND Y = 105 else
"111111111111" when X = 297 AND Y = 105 else
"111111111111" when X = 298 AND Y = 105 else
"111111111111" when X = 299 AND Y = 105 else
"111111111111" when X = 300 AND Y = 105 else
"111111111111" when X = 301 AND Y = 105 else
"111111111111" when X = 302 AND Y = 105 else
"111111111111" when X = 303 AND Y = 105 else
"111111111111" when X = 304 AND Y = 105 else
"110111011111" when X = 305 AND Y = 105 else
"110111011111" when X = 306 AND Y = 105 else
"110111011111" when X = 307 AND Y = 105 else
"110111011111" when X = 308 AND Y = 105 else
"110111011111" when X = 309 AND Y = 105 else
"110111011111" when X = 310 AND Y = 105 else
"110111011111" when X = 311 AND Y = 105 else
"110111011111" when X = 312 AND Y = 105 else
"110111011111" when X = 313 AND Y = 105 else
"110111011111" when X = 314 AND Y = 105 else
"110111011111" when X = 315 AND Y = 105 else
"110111011111" when X = 316 AND Y = 105 else
"110111011111" when X = 317 AND Y = 105 else
"110111011111" when X = 318 AND Y = 105 else
"110111011111" when X = 319 AND Y = 105 else
"110111011111" when X = 320 AND Y = 105 else
"110111011111" when X = 321 AND Y = 105 else
"110111011111" when X = 322 AND Y = 105 else
"110111011111" when X = 323 AND Y = 105 else
"110111011111" when X = 324 AND Y = 105 else
"100010011101" when X = 0 AND Y = 106 else
"100010011101" when X = 1 AND Y = 106 else
"100010011101" when X = 2 AND Y = 106 else
"100010011101" when X = 3 AND Y = 106 else
"100010011101" when X = 4 AND Y = 106 else
"100010011101" when X = 5 AND Y = 106 else
"100010011101" when X = 6 AND Y = 106 else
"100010011101" when X = 7 AND Y = 106 else
"100010011101" when X = 8 AND Y = 106 else
"100010011101" when X = 9 AND Y = 106 else
"100010011101" when X = 10 AND Y = 106 else
"100010011101" when X = 11 AND Y = 106 else
"100010011101" when X = 12 AND Y = 106 else
"100010011101" when X = 13 AND Y = 106 else
"100010011101" when X = 14 AND Y = 106 else
"100010011101" when X = 15 AND Y = 106 else
"100010011101" when X = 16 AND Y = 106 else
"100010011101" when X = 17 AND Y = 106 else
"100010011101" when X = 18 AND Y = 106 else
"100010011101" when X = 19 AND Y = 106 else
"100010011101" when X = 20 AND Y = 106 else
"100010011101" when X = 21 AND Y = 106 else
"100010011101" when X = 22 AND Y = 106 else
"100010011101" when X = 23 AND Y = 106 else
"100010011101" when X = 24 AND Y = 106 else
"110111011111" when X = 25 AND Y = 106 else
"110111011111" when X = 26 AND Y = 106 else
"110111011111" when X = 27 AND Y = 106 else
"110111011111" when X = 28 AND Y = 106 else
"110111011111" when X = 29 AND Y = 106 else
"110111011111" when X = 30 AND Y = 106 else
"110111011111" when X = 31 AND Y = 106 else
"110111011111" when X = 32 AND Y = 106 else
"110111011111" when X = 33 AND Y = 106 else
"110111011111" when X = 34 AND Y = 106 else
"110111011111" when X = 35 AND Y = 106 else
"110111011111" when X = 36 AND Y = 106 else
"110111011111" when X = 37 AND Y = 106 else
"110111011111" when X = 38 AND Y = 106 else
"110111011111" when X = 39 AND Y = 106 else
"110111011111" when X = 40 AND Y = 106 else
"110111011111" when X = 41 AND Y = 106 else
"110111011111" when X = 42 AND Y = 106 else
"110111011111" when X = 43 AND Y = 106 else
"110111011111" when X = 44 AND Y = 106 else
"110111011111" when X = 45 AND Y = 106 else
"110111011111" when X = 46 AND Y = 106 else
"110111011111" when X = 47 AND Y = 106 else
"110111011111" when X = 48 AND Y = 106 else
"110111011111" when X = 49 AND Y = 106 else
"110111011111" when X = 50 AND Y = 106 else
"110111011111" when X = 51 AND Y = 106 else
"110111011111" when X = 52 AND Y = 106 else
"110111011111" when X = 53 AND Y = 106 else
"110111011111" when X = 54 AND Y = 106 else
"110111011111" when X = 55 AND Y = 106 else
"110111011111" when X = 56 AND Y = 106 else
"110111011111" when X = 57 AND Y = 106 else
"110111011111" when X = 58 AND Y = 106 else
"110111011111" when X = 59 AND Y = 106 else
"110111011111" when X = 60 AND Y = 106 else
"110111011111" when X = 61 AND Y = 106 else
"110111011111" when X = 62 AND Y = 106 else
"110111011111" when X = 63 AND Y = 106 else
"110111011111" when X = 64 AND Y = 106 else
"110111011111" when X = 65 AND Y = 106 else
"110111011111" when X = 66 AND Y = 106 else
"110111011111" when X = 67 AND Y = 106 else
"110111011111" when X = 68 AND Y = 106 else
"110111011111" when X = 69 AND Y = 106 else
"111111111111" when X = 70 AND Y = 106 else
"111111111111" when X = 71 AND Y = 106 else
"111111111111" when X = 72 AND Y = 106 else
"111111111111" when X = 73 AND Y = 106 else
"111111111111" when X = 74 AND Y = 106 else
"111111111111" when X = 75 AND Y = 106 else
"111111111111" when X = 76 AND Y = 106 else
"111111111111" when X = 77 AND Y = 106 else
"111111111111" when X = 78 AND Y = 106 else
"111111111111" when X = 79 AND Y = 106 else
"111111111111" when X = 80 AND Y = 106 else
"111111111111" when X = 81 AND Y = 106 else
"111111111111" when X = 82 AND Y = 106 else
"111111111111" when X = 83 AND Y = 106 else
"111111111111" when X = 84 AND Y = 106 else
"111111111111" when X = 85 AND Y = 106 else
"111111111111" when X = 86 AND Y = 106 else
"111111111111" when X = 87 AND Y = 106 else
"111111111111" when X = 88 AND Y = 106 else
"111111111111" when X = 89 AND Y = 106 else
"111111111111" when X = 90 AND Y = 106 else
"111111111111" when X = 91 AND Y = 106 else
"111111111111" when X = 92 AND Y = 106 else
"111111111111" when X = 93 AND Y = 106 else
"111111111111" when X = 94 AND Y = 106 else
"111111111111" when X = 95 AND Y = 106 else
"111111111111" when X = 96 AND Y = 106 else
"111111111111" when X = 97 AND Y = 106 else
"111111111111" when X = 98 AND Y = 106 else
"111111111111" when X = 99 AND Y = 106 else
"111111111111" when X = 100 AND Y = 106 else
"111111111111" when X = 101 AND Y = 106 else
"111111111111" when X = 102 AND Y = 106 else
"111111111111" when X = 103 AND Y = 106 else
"111111111111" when X = 104 AND Y = 106 else
"111111111111" when X = 105 AND Y = 106 else
"111111111111" when X = 106 AND Y = 106 else
"111111111111" when X = 107 AND Y = 106 else
"111111111111" when X = 108 AND Y = 106 else
"111111111111" when X = 109 AND Y = 106 else
"111111111111" when X = 110 AND Y = 106 else
"111111111111" when X = 111 AND Y = 106 else
"111111111111" when X = 112 AND Y = 106 else
"111111111111" when X = 113 AND Y = 106 else
"111111111111" when X = 114 AND Y = 106 else
"111111111111" when X = 115 AND Y = 106 else
"111111111111" when X = 116 AND Y = 106 else
"111111111111" when X = 117 AND Y = 106 else
"111111111111" when X = 118 AND Y = 106 else
"111111111111" when X = 119 AND Y = 106 else
"111111111111" when X = 120 AND Y = 106 else
"111111111111" when X = 121 AND Y = 106 else
"111111111111" when X = 122 AND Y = 106 else
"111111111111" when X = 123 AND Y = 106 else
"111111111111" when X = 124 AND Y = 106 else
"111111111111" when X = 125 AND Y = 106 else
"111111111111" when X = 126 AND Y = 106 else
"111111111111" when X = 127 AND Y = 106 else
"111111111111" when X = 128 AND Y = 106 else
"111111111111" when X = 129 AND Y = 106 else
"111111111111" when X = 130 AND Y = 106 else
"111111111111" when X = 131 AND Y = 106 else
"111111111111" when X = 132 AND Y = 106 else
"111111111111" when X = 133 AND Y = 106 else
"111111111111" when X = 134 AND Y = 106 else
"111111111111" when X = 135 AND Y = 106 else
"111111111111" when X = 136 AND Y = 106 else
"111111111111" when X = 137 AND Y = 106 else
"111111111111" when X = 138 AND Y = 106 else
"111111111111" when X = 139 AND Y = 106 else
"111111111111" when X = 140 AND Y = 106 else
"111111111111" when X = 141 AND Y = 106 else
"111111111111" when X = 142 AND Y = 106 else
"111111111111" when X = 143 AND Y = 106 else
"111111111111" when X = 144 AND Y = 106 else
"111111111111" when X = 145 AND Y = 106 else
"111111111111" when X = 146 AND Y = 106 else
"111111111111" when X = 147 AND Y = 106 else
"111111111111" when X = 148 AND Y = 106 else
"111111111111" when X = 149 AND Y = 106 else
"111111111111" when X = 150 AND Y = 106 else
"111111111111" when X = 151 AND Y = 106 else
"111111111111" when X = 152 AND Y = 106 else
"111111111111" when X = 153 AND Y = 106 else
"111111111111" when X = 154 AND Y = 106 else
"111111111111" when X = 155 AND Y = 106 else
"111111111111" when X = 156 AND Y = 106 else
"111111111111" when X = 157 AND Y = 106 else
"111111111111" when X = 158 AND Y = 106 else
"111111111111" when X = 159 AND Y = 106 else
"110111011111" when X = 160 AND Y = 106 else
"110111011111" when X = 161 AND Y = 106 else
"110111011111" when X = 162 AND Y = 106 else
"110111011111" when X = 163 AND Y = 106 else
"110111011111" when X = 164 AND Y = 106 else
"110111011111" when X = 165 AND Y = 106 else
"110111011111" when X = 166 AND Y = 106 else
"110111011111" when X = 167 AND Y = 106 else
"110111011111" when X = 168 AND Y = 106 else
"110111011111" when X = 169 AND Y = 106 else
"110111011111" when X = 170 AND Y = 106 else
"110111011111" when X = 171 AND Y = 106 else
"110111011111" when X = 172 AND Y = 106 else
"110111011111" when X = 173 AND Y = 106 else
"110111011111" when X = 174 AND Y = 106 else
"110111011111" when X = 175 AND Y = 106 else
"110111011111" when X = 176 AND Y = 106 else
"110111011111" when X = 177 AND Y = 106 else
"110111011111" when X = 178 AND Y = 106 else
"110111011111" when X = 179 AND Y = 106 else
"110111011111" when X = 180 AND Y = 106 else
"110111011111" when X = 181 AND Y = 106 else
"110111011111" when X = 182 AND Y = 106 else
"110111011111" when X = 183 AND Y = 106 else
"110111011111" when X = 184 AND Y = 106 else
"110111011111" when X = 185 AND Y = 106 else
"110111011111" when X = 186 AND Y = 106 else
"110111011111" when X = 187 AND Y = 106 else
"110111011111" when X = 188 AND Y = 106 else
"110111011111" when X = 189 AND Y = 106 else
"110111011111" when X = 190 AND Y = 106 else
"110111011111" when X = 191 AND Y = 106 else
"110111011111" when X = 192 AND Y = 106 else
"110111011111" when X = 193 AND Y = 106 else
"110111011111" when X = 194 AND Y = 106 else
"110111011111" when X = 195 AND Y = 106 else
"110111011111" when X = 196 AND Y = 106 else
"110111011111" when X = 197 AND Y = 106 else
"110111011111" when X = 198 AND Y = 106 else
"110111011111" when X = 199 AND Y = 106 else
"110111011111" when X = 200 AND Y = 106 else
"110111011111" when X = 201 AND Y = 106 else
"110111011111" when X = 202 AND Y = 106 else
"110111011111" when X = 203 AND Y = 106 else
"110111011111" when X = 204 AND Y = 106 else
"111111111111" when X = 205 AND Y = 106 else
"111111111111" when X = 206 AND Y = 106 else
"111111111111" when X = 207 AND Y = 106 else
"111111111111" when X = 208 AND Y = 106 else
"111111111111" when X = 209 AND Y = 106 else
"111111111111" when X = 210 AND Y = 106 else
"111111111111" when X = 211 AND Y = 106 else
"111111111111" when X = 212 AND Y = 106 else
"111111111111" when X = 213 AND Y = 106 else
"111111111111" when X = 214 AND Y = 106 else
"110111011111" when X = 215 AND Y = 106 else
"110111011111" when X = 216 AND Y = 106 else
"110111011111" when X = 217 AND Y = 106 else
"110111011111" when X = 218 AND Y = 106 else
"110111011111" when X = 219 AND Y = 106 else
"110111011111" when X = 220 AND Y = 106 else
"110111011111" when X = 221 AND Y = 106 else
"110111011111" when X = 222 AND Y = 106 else
"110111011111" when X = 223 AND Y = 106 else
"110111011111" when X = 224 AND Y = 106 else
"110111011111" when X = 225 AND Y = 106 else
"110111011111" when X = 226 AND Y = 106 else
"110111011111" when X = 227 AND Y = 106 else
"110111011111" when X = 228 AND Y = 106 else
"110111011111" when X = 229 AND Y = 106 else
"110111011111" when X = 230 AND Y = 106 else
"110111011111" when X = 231 AND Y = 106 else
"110111011111" when X = 232 AND Y = 106 else
"110111011111" when X = 233 AND Y = 106 else
"110111011111" when X = 234 AND Y = 106 else
"110111011111" when X = 235 AND Y = 106 else
"110111011111" when X = 236 AND Y = 106 else
"110111011111" when X = 237 AND Y = 106 else
"110111011111" when X = 238 AND Y = 106 else
"110111011111" when X = 239 AND Y = 106 else
"110111011111" when X = 240 AND Y = 106 else
"110111011111" when X = 241 AND Y = 106 else
"110111011111" when X = 242 AND Y = 106 else
"110111011111" when X = 243 AND Y = 106 else
"110111011111" when X = 244 AND Y = 106 else
"110111011111" when X = 245 AND Y = 106 else
"110111011111" when X = 246 AND Y = 106 else
"110111011111" when X = 247 AND Y = 106 else
"110111011111" when X = 248 AND Y = 106 else
"110111011111" when X = 249 AND Y = 106 else
"110111011111" when X = 250 AND Y = 106 else
"110111011111" when X = 251 AND Y = 106 else
"110111011111" when X = 252 AND Y = 106 else
"110111011111" when X = 253 AND Y = 106 else
"110111011111" when X = 254 AND Y = 106 else
"110111011111" when X = 255 AND Y = 106 else
"110111011111" when X = 256 AND Y = 106 else
"110111011111" when X = 257 AND Y = 106 else
"110111011111" when X = 258 AND Y = 106 else
"110111011111" when X = 259 AND Y = 106 else
"110111011111" when X = 260 AND Y = 106 else
"110111011111" when X = 261 AND Y = 106 else
"110111011111" when X = 262 AND Y = 106 else
"110111011111" when X = 263 AND Y = 106 else
"110111011111" when X = 264 AND Y = 106 else
"110111011111" when X = 265 AND Y = 106 else
"110111011111" when X = 266 AND Y = 106 else
"110111011111" when X = 267 AND Y = 106 else
"110111011111" when X = 268 AND Y = 106 else
"110111011111" when X = 269 AND Y = 106 else
"110111011111" when X = 270 AND Y = 106 else
"110111011111" when X = 271 AND Y = 106 else
"110111011111" when X = 272 AND Y = 106 else
"110111011111" when X = 273 AND Y = 106 else
"110111011111" when X = 274 AND Y = 106 else
"110111011111" when X = 275 AND Y = 106 else
"110111011111" when X = 276 AND Y = 106 else
"110111011111" when X = 277 AND Y = 106 else
"110111011111" when X = 278 AND Y = 106 else
"110111011111" when X = 279 AND Y = 106 else
"111111111111" when X = 280 AND Y = 106 else
"111111111111" when X = 281 AND Y = 106 else
"111111111111" when X = 282 AND Y = 106 else
"111111111111" when X = 283 AND Y = 106 else
"111111111111" when X = 284 AND Y = 106 else
"111111111111" when X = 285 AND Y = 106 else
"111111111111" when X = 286 AND Y = 106 else
"111111111111" when X = 287 AND Y = 106 else
"111111111111" when X = 288 AND Y = 106 else
"111111111111" when X = 289 AND Y = 106 else
"111111111111" when X = 290 AND Y = 106 else
"111111111111" when X = 291 AND Y = 106 else
"111111111111" when X = 292 AND Y = 106 else
"111111111111" when X = 293 AND Y = 106 else
"111111111111" when X = 294 AND Y = 106 else
"111111111111" when X = 295 AND Y = 106 else
"111111111111" when X = 296 AND Y = 106 else
"111111111111" when X = 297 AND Y = 106 else
"111111111111" when X = 298 AND Y = 106 else
"111111111111" when X = 299 AND Y = 106 else
"111111111111" when X = 300 AND Y = 106 else
"111111111111" when X = 301 AND Y = 106 else
"111111111111" when X = 302 AND Y = 106 else
"111111111111" when X = 303 AND Y = 106 else
"111111111111" when X = 304 AND Y = 106 else
"110111011111" when X = 305 AND Y = 106 else
"110111011111" when X = 306 AND Y = 106 else
"110111011111" when X = 307 AND Y = 106 else
"110111011111" when X = 308 AND Y = 106 else
"110111011111" when X = 309 AND Y = 106 else
"110111011111" when X = 310 AND Y = 106 else
"110111011111" when X = 311 AND Y = 106 else
"110111011111" when X = 312 AND Y = 106 else
"110111011111" when X = 313 AND Y = 106 else
"110111011111" when X = 314 AND Y = 106 else
"110111011111" when X = 315 AND Y = 106 else
"110111011111" when X = 316 AND Y = 106 else
"110111011111" when X = 317 AND Y = 106 else
"110111011111" when X = 318 AND Y = 106 else
"110111011111" when X = 319 AND Y = 106 else
"110111011111" when X = 320 AND Y = 106 else
"110111011111" when X = 321 AND Y = 106 else
"110111011111" when X = 322 AND Y = 106 else
"110111011111" when X = 323 AND Y = 106 else
"110111011111" when X = 324 AND Y = 106 else
"100010011101" when X = 0 AND Y = 107 else
"100010011101" when X = 1 AND Y = 107 else
"100010011101" when X = 2 AND Y = 107 else
"100010011101" when X = 3 AND Y = 107 else
"100010011101" when X = 4 AND Y = 107 else
"100010011101" when X = 5 AND Y = 107 else
"100010011101" when X = 6 AND Y = 107 else
"100010011101" when X = 7 AND Y = 107 else
"100010011101" when X = 8 AND Y = 107 else
"100010011101" when X = 9 AND Y = 107 else
"100010011101" when X = 10 AND Y = 107 else
"100010011101" when X = 11 AND Y = 107 else
"100010011101" when X = 12 AND Y = 107 else
"100010011101" when X = 13 AND Y = 107 else
"100010011101" when X = 14 AND Y = 107 else
"100010011101" when X = 15 AND Y = 107 else
"100010011101" when X = 16 AND Y = 107 else
"100010011101" when X = 17 AND Y = 107 else
"100010011101" when X = 18 AND Y = 107 else
"100010011101" when X = 19 AND Y = 107 else
"100010011101" when X = 20 AND Y = 107 else
"100010011101" when X = 21 AND Y = 107 else
"100010011101" when X = 22 AND Y = 107 else
"100010011101" when X = 23 AND Y = 107 else
"100010011101" when X = 24 AND Y = 107 else
"110111011111" when X = 25 AND Y = 107 else
"110111011111" when X = 26 AND Y = 107 else
"110111011111" when X = 27 AND Y = 107 else
"110111011111" when X = 28 AND Y = 107 else
"110111011111" when X = 29 AND Y = 107 else
"110111011111" when X = 30 AND Y = 107 else
"110111011111" when X = 31 AND Y = 107 else
"110111011111" when X = 32 AND Y = 107 else
"110111011111" when X = 33 AND Y = 107 else
"110111011111" when X = 34 AND Y = 107 else
"110111011111" when X = 35 AND Y = 107 else
"110111011111" when X = 36 AND Y = 107 else
"110111011111" when X = 37 AND Y = 107 else
"110111011111" when X = 38 AND Y = 107 else
"110111011111" when X = 39 AND Y = 107 else
"110111011111" when X = 40 AND Y = 107 else
"110111011111" when X = 41 AND Y = 107 else
"110111011111" when X = 42 AND Y = 107 else
"110111011111" when X = 43 AND Y = 107 else
"110111011111" when X = 44 AND Y = 107 else
"110111011111" when X = 45 AND Y = 107 else
"110111011111" when X = 46 AND Y = 107 else
"110111011111" when X = 47 AND Y = 107 else
"110111011111" when X = 48 AND Y = 107 else
"110111011111" when X = 49 AND Y = 107 else
"110111011111" when X = 50 AND Y = 107 else
"110111011111" when X = 51 AND Y = 107 else
"110111011111" when X = 52 AND Y = 107 else
"110111011111" when X = 53 AND Y = 107 else
"110111011111" when X = 54 AND Y = 107 else
"110111011111" when X = 55 AND Y = 107 else
"110111011111" when X = 56 AND Y = 107 else
"110111011111" when X = 57 AND Y = 107 else
"110111011111" when X = 58 AND Y = 107 else
"110111011111" when X = 59 AND Y = 107 else
"110111011111" when X = 60 AND Y = 107 else
"110111011111" when X = 61 AND Y = 107 else
"110111011111" when X = 62 AND Y = 107 else
"110111011111" when X = 63 AND Y = 107 else
"110111011111" when X = 64 AND Y = 107 else
"110111011111" when X = 65 AND Y = 107 else
"110111011111" when X = 66 AND Y = 107 else
"110111011111" when X = 67 AND Y = 107 else
"110111011111" when X = 68 AND Y = 107 else
"110111011111" when X = 69 AND Y = 107 else
"111111111111" when X = 70 AND Y = 107 else
"111111111111" when X = 71 AND Y = 107 else
"111111111111" when X = 72 AND Y = 107 else
"111111111111" when X = 73 AND Y = 107 else
"111111111111" when X = 74 AND Y = 107 else
"111111111111" when X = 75 AND Y = 107 else
"111111111111" when X = 76 AND Y = 107 else
"111111111111" when X = 77 AND Y = 107 else
"111111111111" when X = 78 AND Y = 107 else
"111111111111" when X = 79 AND Y = 107 else
"111111111111" when X = 80 AND Y = 107 else
"111111111111" when X = 81 AND Y = 107 else
"111111111111" when X = 82 AND Y = 107 else
"111111111111" when X = 83 AND Y = 107 else
"111111111111" when X = 84 AND Y = 107 else
"111111111111" when X = 85 AND Y = 107 else
"111111111111" when X = 86 AND Y = 107 else
"111111111111" when X = 87 AND Y = 107 else
"111111111111" when X = 88 AND Y = 107 else
"111111111111" when X = 89 AND Y = 107 else
"111111111111" when X = 90 AND Y = 107 else
"111111111111" when X = 91 AND Y = 107 else
"111111111111" when X = 92 AND Y = 107 else
"111111111111" when X = 93 AND Y = 107 else
"111111111111" when X = 94 AND Y = 107 else
"111111111111" when X = 95 AND Y = 107 else
"111111111111" when X = 96 AND Y = 107 else
"111111111111" when X = 97 AND Y = 107 else
"111111111111" when X = 98 AND Y = 107 else
"111111111111" when X = 99 AND Y = 107 else
"111111111111" when X = 100 AND Y = 107 else
"111111111111" when X = 101 AND Y = 107 else
"111111111111" when X = 102 AND Y = 107 else
"111111111111" when X = 103 AND Y = 107 else
"111111111111" when X = 104 AND Y = 107 else
"111111111111" when X = 105 AND Y = 107 else
"111111111111" when X = 106 AND Y = 107 else
"111111111111" when X = 107 AND Y = 107 else
"111111111111" when X = 108 AND Y = 107 else
"111111111111" when X = 109 AND Y = 107 else
"111111111111" when X = 110 AND Y = 107 else
"111111111111" when X = 111 AND Y = 107 else
"111111111111" when X = 112 AND Y = 107 else
"111111111111" when X = 113 AND Y = 107 else
"111111111111" when X = 114 AND Y = 107 else
"111111111111" when X = 115 AND Y = 107 else
"111111111111" when X = 116 AND Y = 107 else
"111111111111" when X = 117 AND Y = 107 else
"111111111111" when X = 118 AND Y = 107 else
"111111111111" when X = 119 AND Y = 107 else
"111111111111" when X = 120 AND Y = 107 else
"111111111111" when X = 121 AND Y = 107 else
"111111111111" when X = 122 AND Y = 107 else
"111111111111" when X = 123 AND Y = 107 else
"111111111111" when X = 124 AND Y = 107 else
"111111111111" when X = 125 AND Y = 107 else
"111111111111" when X = 126 AND Y = 107 else
"111111111111" when X = 127 AND Y = 107 else
"111111111111" when X = 128 AND Y = 107 else
"111111111111" when X = 129 AND Y = 107 else
"111111111111" when X = 130 AND Y = 107 else
"111111111111" when X = 131 AND Y = 107 else
"111111111111" when X = 132 AND Y = 107 else
"111111111111" when X = 133 AND Y = 107 else
"111111111111" when X = 134 AND Y = 107 else
"111111111111" when X = 135 AND Y = 107 else
"111111111111" when X = 136 AND Y = 107 else
"111111111111" when X = 137 AND Y = 107 else
"111111111111" when X = 138 AND Y = 107 else
"111111111111" when X = 139 AND Y = 107 else
"111111111111" when X = 140 AND Y = 107 else
"111111111111" when X = 141 AND Y = 107 else
"111111111111" when X = 142 AND Y = 107 else
"111111111111" when X = 143 AND Y = 107 else
"111111111111" when X = 144 AND Y = 107 else
"111111111111" when X = 145 AND Y = 107 else
"111111111111" when X = 146 AND Y = 107 else
"111111111111" when X = 147 AND Y = 107 else
"111111111111" when X = 148 AND Y = 107 else
"111111111111" when X = 149 AND Y = 107 else
"111111111111" when X = 150 AND Y = 107 else
"111111111111" when X = 151 AND Y = 107 else
"111111111111" when X = 152 AND Y = 107 else
"111111111111" when X = 153 AND Y = 107 else
"111111111111" when X = 154 AND Y = 107 else
"111111111111" when X = 155 AND Y = 107 else
"111111111111" when X = 156 AND Y = 107 else
"111111111111" when X = 157 AND Y = 107 else
"111111111111" when X = 158 AND Y = 107 else
"111111111111" when X = 159 AND Y = 107 else
"110111011111" when X = 160 AND Y = 107 else
"110111011111" when X = 161 AND Y = 107 else
"110111011111" when X = 162 AND Y = 107 else
"110111011111" when X = 163 AND Y = 107 else
"110111011111" when X = 164 AND Y = 107 else
"110111011111" when X = 165 AND Y = 107 else
"110111011111" when X = 166 AND Y = 107 else
"110111011111" when X = 167 AND Y = 107 else
"110111011111" when X = 168 AND Y = 107 else
"110111011111" when X = 169 AND Y = 107 else
"110111011111" when X = 170 AND Y = 107 else
"110111011111" when X = 171 AND Y = 107 else
"110111011111" when X = 172 AND Y = 107 else
"110111011111" when X = 173 AND Y = 107 else
"110111011111" when X = 174 AND Y = 107 else
"110111011111" when X = 175 AND Y = 107 else
"110111011111" when X = 176 AND Y = 107 else
"110111011111" when X = 177 AND Y = 107 else
"110111011111" when X = 178 AND Y = 107 else
"110111011111" when X = 179 AND Y = 107 else
"110111011111" when X = 180 AND Y = 107 else
"110111011111" when X = 181 AND Y = 107 else
"110111011111" when X = 182 AND Y = 107 else
"110111011111" when X = 183 AND Y = 107 else
"110111011111" when X = 184 AND Y = 107 else
"110111011111" when X = 185 AND Y = 107 else
"110111011111" when X = 186 AND Y = 107 else
"110111011111" when X = 187 AND Y = 107 else
"110111011111" when X = 188 AND Y = 107 else
"110111011111" when X = 189 AND Y = 107 else
"110111011111" when X = 190 AND Y = 107 else
"110111011111" when X = 191 AND Y = 107 else
"110111011111" when X = 192 AND Y = 107 else
"110111011111" when X = 193 AND Y = 107 else
"110111011111" when X = 194 AND Y = 107 else
"110111011111" when X = 195 AND Y = 107 else
"110111011111" when X = 196 AND Y = 107 else
"110111011111" when X = 197 AND Y = 107 else
"110111011111" when X = 198 AND Y = 107 else
"110111011111" when X = 199 AND Y = 107 else
"110111011111" when X = 200 AND Y = 107 else
"110111011111" when X = 201 AND Y = 107 else
"110111011111" when X = 202 AND Y = 107 else
"110111011111" when X = 203 AND Y = 107 else
"110111011111" when X = 204 AND Y = 107 else
"111111111111" when X = 205 AND Y = 107 else
"111111111111" when X = 206 AND Y = 107 else
"111111111111" when X = 207 AND Y = 107 else
"111111111111" when X = 208 AND Y = 107 else
"111111111111" when X = 209 AND Y = 107 else
"111111111111" when X = 210 AND Y = 107 else
"111111111111" when X = 211 AND Y = 107 else
"111111111111" when X = 212 AND Y = 107 else
"111111111111" when X = 213 AND Y = 107 else
"111111111111" when X = 214 AND Y = 107 else
"110111011111" when X = 215 AND Y = 107 else
"110111011111" when X = 216 AND Y = 107 else
"110111011111" when X = 217 AND Y = 107 else
"110111011111" when X = 218 AND Y = 107 else
"110111011111" when X = 219 AND Y = 107 else
"110111011111" when X = 220 AND Y = 107 else
"110111011111" when X = 221 AND Y = 107 else
"110111011111" when X = 222 AND Y = 107 else
"110111011111" when X = 223 AND Y = 107 else
"110111011111" when X = 224 AND Y = 107 else
"110111011111" when X = 225 AND Y = 107 else
"110111011111" when X = 226 AND Y = 107 else
"110111011111" when X = 227 AND Y = 107 else
"110111011111" when X = 228 AND Y = 107 else
"110111011111" when X = 229 AND Y = 107 else
"110111011111" when X = 230 AND Y = 107 else
"110111011111" when X = 231 AND Y = 107 else
"110111011111" when X = 232 AND Y = 107 else
"110111011111" when X = 233 AND Y = 107 else
"110111011111" when X = 234 AND Y = 107 else
"110111011111" when X = 235 AND Y = 107 else
"110111011111" when X = 236 AND Y = 107 else
"110111011111" when X = 237 AND Y = 107 else
"110111011111" when X = 238 AND Y = 107 else
"110111011111" when X = 239 AND Y = 107 else
"110111011111" when X = 240 AND Y = 107 else
"110111011111" when X = 241 AND Y = 107 else
"110111011111" when X = 242 AND Y = 107 else
"110111011111" when X = 243 AND Y = 107 else
"110111011111" when X = 244 AND Y = 107 else
"110111011111" when X = 245 AND Y = 107 else
"110111011111" when X = 246 AND Y = 107 else
"110111011111" when X = 247 AND Y = 107 else
"110111011111" when X = 248 AND Y = 107 else
"110111011111" when X = 249 AND Y = 107 else
"110111011111" when X = 250 AND Y = 107 else
"110111011111" when X = 251 AND Y = 107 else
"110111011111" when X = 252 AND Y = 107 else
"110111011111" when X = 253 AND Y = 107 else
"110111011111" when X = 254 AND Y = 107 else
"110111011111" when X = 255 AND Y = 107 else
"110111011111" when X = 256 AND Y = 107 else
"110111011111" when X = 257 AND Y = 107 else
"110111011111" when X = 258 AND Y = 107 else
"110111011111" when X = 259 AND Y = 107 else
"110111011111" when X = 260 AND Y = 107 else
"110111011111" when X = 261 AND Y = 107 else
"110111011111" when X = 262 AND Y = 107 else
"110111011111" when X = 263 AND Y = 107 else
"110111011111" when X = 264 AND Y = 107 else
"110111011111" when X = 265 AND Y = 107 else
"110111011111" when X = 266 AND Y = 107 else
"110111011111" when X = 267 AND Y = 107 else
"110111011111" when X = 268 AND Y = 107 else
"110111011111" when X = 269 AND Y = 107 else
"110111011111" when X = 270 AND Y = 107 else
"110111011111" when X = 271 AND Y = 107 else
"110111011111" when X = 272 AND Y = 107 else
"110111011111" when X = 273 AND Y = 107 else
"110111011111" when X = 274 AND Y = 107 else
"110111011111" when X = 275 AND Y = 107 else
"110111011111" when X = 276 AND Y = 107 else
"110111011111" when X = 277 AND Y = 107 else
"110111011111" when X = 278 AND Y = 107 else
"110111011111" when X = 279 AND Y = 107 else
"111111111111" when X = 280 AND Y = 107 else
"111111111111" when X = 281 AND Y = 107 else
"111111111111" when X = 282 AND Y = 107 else
"111111111111" when X = 283 AND Y = 107 else
"111111111111" when X = 284 AND Y = 107 else
"111111111111" when X = 285 AND Y = 107 else
"111111111111" when X = 286 AND Y = 107 else
"111111111111" when X = 287 AND Y = 107 else
"111111111111" when X = 288 AND Y = 107 else
"111111111111" when X = 289 AND Y = 107 else
"111111111111" when X = 290 AND Y = 107 else
"111111111111" when X = 291 AND Y = 107 else
"111111111111" when X = 292 AND Y = 107 else
"111111111111" when X = 293 AND Y = 107 else
"111111111111" when X = 294 AND Y = 107 else
"111111111111" when X = 295 AND Y = 107 else
"111111111111" when X = 296 AND Y = 107 else
"111111111111" when X = 297 AND Y = 107 else
"111111111111" when X = 298 AND Y = 107 else
"111111111111" when X = 299 AND Y = 107 else
"111111111111" when X = 300 AND Y = 107 else
"111111111111" when X = 301 AND Y = 107 else
"111111111111" when X = 302 AND Y = 107 else
"111111111111" when X = 303 AND Y = 107 else
"111111111111" when X = 304 AND Y = 107 else
"110111011111" when X = 305 AND Y = 107 else
"110111011111" when X = 306 AND Y = 107 else
"110111011111" when X = 307 AND Y = 107 else
"110111011111" when X = 308 AND Y = 107 else
"110111011111" when X = 309 AND Y = 107 else
"110111011111" when X = 310 AND Y = 107 else
"110111011111" when X = 311 AND Y = 107 else
"110111011111" when X = 312 AND Y = 107 else
"110111011111" when X = 313 AND Y = 107 else
"110111011111" when X = 314 AND Y = 107 else
"110111011111" when X = 315 AND Y = 107 else
"110111011111" when X = 316 AND Y = 107 else
"110111011111" when X = 317 AND Y = 107 else
"110111011111" when X = 318 AND Y = 107 else
"110111011111" when X = 319 AND Y = 107 else
"110111011111" when X = 320 AND Y = 107 else
"110111011111" when X = 321 AND Y = 107 else
"110111011111" when X = 322 AND Y = 107 else
"110111011111" when X = 323 AND Y = 107 else
"110111011111" when X = 324 AND Y = 107 else
"100010011101" when X = 0 AND Y = 108 else
"100010011101" when X = 1 AND Y = 108 else
"100010011101" when X = 2 AND Y = 108 else
"100010011101" when X = 3 AND Y = 108 else
"100010011101" when X = 4 AND Y = 108 else
"100010011101" when X = 5 AND Y = 108 else
"100010011101" when X = 6 AND Y = 108 else
"100010011101" when X = 7 AND Y = 108 else
"100010011101" when X = 8 AND Y = 108 else
"100010011101" when X = 9 AND Y = 108 else
"100010011101" when X = 10 AND Y = 108 else
"100010011101" when X = 11 AND Y = 108 else
"100010011101" when X = 12 AND Y = 108 else
"100010011101" when X = 13 AND Y = 108 else
"100010011101" when X = 14 AND Y = 108 else
"100010011101" when X = 15 AND Y = 108 else
"100010011101" when X = 16 AND Y = 108 else
"100010011101" when X = 17 AND Y = 108 else
"100010011101" when X = 18 AND Y = 108 else
"100010011101" when X = 19 AND Y = 108 else
"100010011101" when X = 20 AND Y = 108 else
"100010011101" when X = 21 AND Y = 108 else
"100010011101" when X = 22 AND Y = 108 else
"100010011101" when X = 23 AND Y = 108 else
"100010011101" when X = 24 AND Y = 108 else
"110111011111" when X = 25 AND Y = 108 else
"110111011111" when X = 26 AND Y = 108 else
"110111011111" when X = 27 AND Y = 108 else
"110111011111" when X = 28 AND Y = 108 else
"110111011111" when X = 29 AND Y = 108 else
"110111011111" when X = 30 AND Y = 108 else
"110111011111" when X = 31 AND Y = 108 else
"110111011111" when X = 32 AND Y = 108 else
"110111011111" when X = 33 AND Y = 108 else
"110111011111" when X = 34 AND Y = 108 else
"110111011111" when X = 35 AND Y = 108 else
"110111011111" when X = 36 AND Y = 108 else
"110111011111" when X = 37 AND Y = 108 else
"110111011111" when X = 38 AND Y = 108 else
"110111011111" when X = 39 AND Y = 108 else
"110111011111" when X = 40 AND Y = 108 else
"110111011111" when X = 41 AND Y = 108 else
"110111011111" when X = 42 AND Y = 108 else
"110111011111" when X = 43 AND Y = 108 else
"110111011111" when X = 44 AND Y = 108 else
"110111011111" when X = 45 AND Y = 108 else
"110111011111" when X = 46 AND Y = 108 else
"110111011111" when X = 47 AND Y = 108 else
"110111011111" when X = 48 AND Y = 108 else
"110111011111" when X = 49 AND Y = 108 else
"110111011111" when X = 50 AND Y = 108 else
"110111011111" when X = 51 AND Y = 108 else
"110111011111" when X = 52 AND Y = 108 else
"110111011111" when X = 53 AND Y = 108 else
"110111011111" when X = 54 AND Y = 108 else
"110111011111" when X = 55 AND Y = 108 else
"110111011111" when X = 56 AND Y = 108 else
"110111011111" when X = 57 AND Y = 108 else
"110111011111" when X = 58 AND Y = 108 else
"110111011111" when X = 59 AND Y = 108 else
"110111011111" when X = 60 AND Y = 108 else
"110111011111" when X = 61 AND Y = 108 else
"110111011111" when X = 62 AND Y = 108 else
"110111011111" when X = 63 AND Y = 108 else
"110111011111" when X = 64 AND Y = 108 else
"110111011111" when X = 65 AND Y = 108 else
"110111011111" when X = 66 AND Y = 108 else
"110111011111" when X = 67 AND Y = 108 else
"110111011111" when X = 68 AND Y = 108 else
"110111011111" when X = 69 AND Y = 108 else
"111111111111" when X = 70 AND Y = 108 else
"111111111111" when X = 71 AND Y = 108 else
"111111111111" when X = 72 AND Y = 108 else
"111111111111" when X = 73 AND Y = 108 else
"111111111111" when X = 74 AND Y = 108 else
"111111111111" when X = 75 AND Y = 108 else
"111111111111" when X = 76 AND Y = 108 else
"111111111111" when X = 77 AND Y = 108 else
"111111111111" when X = 78 AND Y = 108 else
"111111111111" when X = 79 AND Y = 108 else
"111111111111" when X = 80 AND Y = 108 else
"111111111111" when X = 81 AND Y = 108 else
"111111111111" when X = 82 AND Y = 108 else
"111111111111" when X = 83 AND Y = 108 else
"111111111111" when X = 84 AND Y = 108 else
"111111111111" when X = 85 AND Y = 108 else
"111111111111" when X = 86 AND Y = 108 else
"111111111111" when X = 87 AND Y = 108 else
"111111111111" when X = 88 AND Y = 108 else
"111111111111" when X = 89 AND Y = 108 else
"111111111111" when X = 90 AND Y = 108 else
"111111111111" when X = 91 AND Y = 108 else
"111111111111" when X = 92 AND Y = 108 else
"111111111111" when X = 93 AND Y = 108 else
"111111111111" when X = 94 AND Y = 108 else
"111111111111" when X = 95 AND Y = 108 else
"111111111111" when X = 96 AND Y = 108 else
"111111111111" when X = 97 AND Y = 108 else
"111111111111" when X = 98 AND Y = 108 else
"111111111111" when X = 99 AND Y = 108 else
"111111111111" when X = 100 AND Y = 108 else
"111111111111" when X = 101 AND Y = 108 else
"111111111111" when X = 102 AND Y = 108 else
"111111111111" when X = 103 AND Y = 108 else
"111111111111" when X = 104 AND Y = 108 else
"111111111111" when X = 105 AND Y = 108 else
"111111111111" when X = 106 AND Y = 108 else
"111111111111" when X = 107 AND Y = 108 else
"111111111111" when X = 108 AND Y = 108 else
"111111111111" when X = 109 AND Y = 108 else
"111111111111" when X = 110 AND Y = 108 else
"111111111111" when X = 111 AND Y = 108 else
"111111111111" when X = 112 AND Y = 108 else
"111111111111" when X = 113 AND Y = 108 else
"111111111111" when X = 114 AND Y = 108 else
"111111111111" when X = 115 AND Y = 108 else
"111111111111" when X = 116 AND Y = 108 else
"111111111111" when X = 117 AND Y = 108 else
"111111111111" when X = 118 AND Y = 108 else
"111111111111" when X = 119 AND Y = 108 else
"111111111111" when X = 120 AND Y = 108 else
"111111111111" when X = 121 AND Y = 108 else
"111111111111" when X = 122 AND Y = 108 else
"111111111111" when X = 123 AND Y = 108 else
"111111111111" when X = 124 AND Y = 108 else
"111111111111" when X = 125 AND Y = 108 else
"111111111111" when X = 126 AND Y = 108 else
"111111111111" when X = 127 AND Y = 108 else
"111111111111" when X = 128 AND Y = 108 else
"111111111111" when X = 129 AND Y = 108 else
"111111111111" when X = 130 AND Y = 108 else
"111111111111" when X = 131 AND Y = 108 else
"111111111111" when X = 132 AND Y = 108 else
"111111111111" when X = 133 AND Y = 108 else
"111111111111" when X = 134 AND Y = 108 else
"111111111111" when X = 135 AND Y = 108 else
"111111111111" when X = 136 AND Y = 108 else
"111111111111" when X = 137 AND Y = 108 else
"111111111111" when X = 138 AND Y = 108 else
"111111111111" when X = 139 AND Y = 108 else
"111111111111" when X = 140 AND Y = 108 else
"111111111111" when X = 141 AND Y = 108 else
"111111111111" when X = 142 AND Y = 108 else
"111111111111" when X = 143 AND Y = 108 else
"111111111111" when X = 144 AND Y = 108 else
"111111111111" when X = 145 AND Y = 108 else
"111111111111" when X = 146 AND Y = 108 else
"111111111111" when X = 147 AND Y = 108 else
"111111111111" when X = 148 AND Y = 108 else
"111111111111" when X = 149 AND Y = 108 else
"111111111111" when X = 150 AND Y = 108 else
"111111111111" when X = 151 AND Y = 108 else
"111111111111" when X = 152 AND Y = 108 else
"111111111111" when X = 153 AND Y = 108 else
"111111111111" when X = 154 AND Y = 108 else
"111111111111" when X = 155 AND Y = 108 else
"111111111111" when X = 156 AND Y = 108 else
"111111111111" when X = 157 AND Y = 108 else
"111111111111" when X = 158 AND Y = 108 else
"111111111111" when X = 159 AND Y = 108 else
"110111011111" when X = 160 AND Y = 108 else
"110111011111" when X = 161 AND Y = 108 else
"110111011111" when X = 162 AND Y = 108 else
"110111011111" when X = 163 AND Y = 108 else
"110111011111" when X = 164 AND Y = 108 else
"110111011111" when X = 165 AND Y = 108 else
"110111011111" when X = 166 AND Y = 108 else
"110111011111" when X = 167 AND Y = 108 else
"110111011111" when X = 168 AND Y = 108 else
"110111011111" when X = 169 AND Y = 108 else
"110111011111" when X = 170 AND Y = 108 else
"110111011111" when X = 171 AND Y = 108 else
"110111011111" when X = 172 AND Y = 108 else
"110111011111" when X = 173 AND Y = 108 else
"110111011111" when X = 174 AND Y = 108 else
"110111011111" when X = 175 AND Y = 108 else
"110111011111" when X = 176 AND Y = 108 else
"110111011111" when X = 177 AND Y = 108 else
"110111011111" when X = 178 AND Y = 108 else
"110111011111" when X = 179 AND Y = 108 else
"110111011111" when X = 180 AND Y = 108 else
"110111011111" when X = 181 AND Y = 108 else
"110111011111" when X = 182 AND Y = 108 else
"110111011111" when X = 183 AND Y = 108 else
"110111011111" when X = 184 AND Y = 108 else
"110111011111" when X = 185 AND Y = 108 else
"110111011111" when X = 186 AND Y = 108 else
"110111011111" when X = 187 AND Y = 108 else
"110111011111" when X = 188 AND Y = 108 else
"110111011111" when X = 189 AND Y = 108 else
"110111011111" when X = 190 AND Y = 108 else
"110111011111" when X = 191 AND Y = 108 else
"110111011111" when X = 192 AND Y = 108 else
"110111011111" when X = 193 AND Y = 108 else
"110111011111" when X = 194 AND Y = 108 else
"110111011111" when X = 195 AND Y = 108 else
"110111011111" when X = 196 AND Y = 108 else
"110111011111" when X = 197 AND Y = 108 else
"110111011111" when X = 198 AND Y = 108 else
"110111011111" when X = 199 AND Y = 108 else
"110111011111" when X = 200 AND Y = 108 else
"110111011111" when X = 201 AND Y = 108 else
"110111011111" when X = 202 AND Y = 108 else
"110111011111" when X = 203 AND Y = 108 else
"110111011111" when X = 204 AND Y = 108 else
"111111111111" when X = 205 AND Y = 108 else
"111111111111" when X = 206 AND Y = 108 else
"111111111111" when X = 207 AND Y = 108 else
"111111111111" when X = 208 AND Y = 108 else
"111111111111" when X = 209 AND Y = 108 else
"111111111111" when X = 210 AND Y = 108 else
"111111111111" when X = 211 AND Y = 108 else
"111111111111" when X = 212 AND Y = 108 else
"111111111111" when X = 213 AND Y = 108 else
"111111111111" when X = 214 AND Y = 108 else
"110111011111" when X = 215 AND Y = 108 else
"110111011111" when X = 216 AND Y = 108 else
"110111011111" when X = 217 AND Y = 108 else
"110111011111" when X = 218 AND Y = 108 else
"110111011111" when X = 219 AND Y = 108 else
"110111011111" when X = 220 AND Y = 108 else
"110111011111" when X = 221 AND Y = 108 else
"110111011111" when X = 222 AND Y = 108 else
"110111011111" when X = 223 AND Y = 108 else
"110111011111" when X = 224 AND Y = 108 else
"110111011111" when X = 225 AND Y = 108 else
"110111011111" when X = 226 AND Y = 108 else
"110111011111" when X = 227 AND Y = 108 else
"110111011111" when X = 228 AND Y = 108 else
"110111011111" when X = 229 AND Y = 108 else
"110111011111" when X = 230 AND Y = 108 else
"110111011111" when X = 231 AND Y = 108 else
"110111011111" when X = 232 AND Y = 108 else
"110111011111" when X = 233 AND Y = 108 else
"110111011111" when X = 234 AND Y = 108 else
"110111011111" when X = 235 AND Y = 108 else
"110111011111" when X = 236 AND Y = 108 else
"110111011111" when X = 237 AND Y = 108 else
"110111011111" when X = 238 AND Y = 108 else
"110111011111" when X = 239 AND Y = 108 else
"110111011111" when X = 240 AND Y = 108 else
"110111011111" when X = 241 AND Y = 108 else
"110111011111" when X = 242 AND Y = 108 else
"110111011111" when X = 243 AND Y = 108 else
"110111011111" when X = 244 AND Y = 108 else
"110111011111" when X = 245 AND Y = 108 else
"110111011111" when X = 246 AND Y = 108 else
"110111011111" when X = 247 AND Y = 108 else
"110111011111" when X = 248 AND Y = 108 else
"110111011111" when X = 249 AND Y = 108 else
"110111011111" when X = 250 AND Y = 108 else
"110111011111" when X = 251 AND Y = 108 else
"110111011111" when X = 252 AND Y = 108 else
"110111011111" when X = 253 AND Y = 108 else
"110111011111" when X = 254 AND Y = 108 else
"110111011111" when X = 255 AND Y = 108 else
"110111011111" when X = 256 AND Y = 108 else
"110111011111" when X = 257 AND Y = 108 else
"110111011111" when X = 258 AND Y = 108 else
"110111011111" when X = 259 AND Y = 108 else
"110111011111" when X = 260 AND Y = 108 else
"110111011111" when X = 261 AND Y = 108 else
"110111011111" when X = 262 AND Y = 108 else
"110111011111" when X = 263 AND Y = 108 else
"110111011111" when X = 264 AND Y = 108 else
"110111011111" when X = 265 AND Y = 108 else
"110111011111" when X = 266 AND Y = 108 else
"110111011111" when X = 267 AND Y = 108 else
"110111011111" when X = 268 AND Y = 108 else
"110111011111" when X = 269 AND Y = 108 else
"110111011111" when X = 270 AND Y = 108 else
"110111011111" when X = 271 AND Y = 108 else
"110111011111" when X = 272 AND Y = 108 else
"110111011111" when X = 273 AND Y = 108 else
"110111011111" when X = 274 AND Y = 108 else
"110111011111" when X = 275 AND Y = 108 else
"110111011111" when X = 276 AND Y = 108 else
"110111011111" when X = 277 AND Y = 108 else
"110111011111" when X = 278 AND Y = 108 else
"110111011111" when X = 279 AND Y = 108 else
"111111111111" when X = 280 AND Y = 108 else
"111111111111" when X = 281 AND Y = 108 else
"111111111111" when X = 282 AND Y = 108 else
"111111111111" when X = 283 AND Y = 108 else
"111111111111" when X = 284 AND Y = 108 else
"111111111111" when X = 285 AND Y = 108 else
"111111111111" when X = 286 AND Y = 108 else
"111111111111" when X = 287 AND Y = 108 else
"111111111111" when X = 288 AND Y = 108 else
"111111111111" when X = 289 AND Y = 108 else
"111111111111" when X = 290 AND Y = 108 else
"111111111111" when X = 291 AND Y = 108 else
"111111111111" when X = 292 AND Y = 108 else
"111111111111" when X = 293 AND Y = 108 else
"111111111111" when X = 294 AND Y = 108 else
"111111111111" when X = 295 AND Y = 108 else
"111111111111" when X = 296 AND Y = 108 else
"111111111111" when X = 297 AND Y = 108 else
"111111111111" when X = 298 AND Y = 108 else
"111111111111" when X = 299 AND Y = 108 else
"111111111111" when X = 300 AND Y = 108 else
"111111111111" when X = 301 AND Y = 108 else
"111111111111" when X = 302 AND Y = 108 else
"111111111111" when X = 303 AND Y = 108 else
"111111111111" when X = 304 AND Y = 108 else
"110111011111" when X = 305 AND Y = 108 else
"110111011111" when X = 306 AND Y = 108 else
"110111011111" when X = 307 AND Y = 108 else
"110111011111" when X = 308 AND Y = 108 else
"110111011111" when X = 309 AND Y = 108 else
"110111011111" when X = 310 AND Y = 108 else
"110111011111" when X = 311 AND Y = 108 else
"110111011111" when X = 312 AND Y = 108 else
"110111011111" when X = 313 AND Y = 108 else
"110111011111" when X = 314 AND Y = 108 else
"110111011111" when X = 315 AND Y = 108 else
"110111011111" when X = 316 AND Y = 108 else
"110111011111" when X = 317 AND Y = 108 else
"110111011111" when X = 318 AND Y = 108 else
"110111011111" when X = 319 AND Y = 108 else
"110111011111" when X = 320 AND Y = 108 else
"110111011111" when X = 321 AND Y = 108 else
"110111011111" when X = 322 AND Y = 108 else
"110111011111" when X = 323 AND Y = 108 else
"110111011111" when X = 324 AND Y = 108 else
"100010011101" when X = 0 AND Y = 109 else
"100010011101" when X = 1 AND Y = 109 else
"100010011101" when X = 2 AND Y = 109 else
"100010011101" when X = 3 AND Y = 109 else
"100010011101" when X = 4 AND Y = 109 else
"100010011101" when X = 5 AND Y = 109 else
"100010011101" when X = 6 AND Y = 109 else
"100010011101" when X = 7 AND Y = 109 else
"100010011101" when X = 8 AND Y = 109 else
"100010011101" when X = 9 AND Y = 109 else
"100010011101" when X = 10 AND Y = 109 else
"100010011101" when X = 11 AND Y = 109 else
"100010011101" when X = 12 AND Y = 109 else
"100010011101" when X = 13 AND Y = 109 else
"100010011101" when X = 14 AND Y = 109 else
"100010011101" when X = 15 AND Y = 109 else
"100010011101" when X = 16 AND Y = 109 else
"100010011101" when X = 17 AND Y = 109 else
"100010011101" when X = 18 AND Y = 109 else
"100010011101" when X = 19 AND Y = 109 else
"100010011101" when X = 20 AND Y = 109 else
"100010011101" when X = 21 AND Y = 109 else
"100010011101" when X = 22 AND Y = 109 else
"100010011101" when X = 23 AND Y = 109 else
"100010011101" when X = 24 AND Y = 109 else
"110111011111" when X = 25 AND Y = 109 else
"110111011111" when X = 26 AND Y = 109 else
"110111011111" when X = 27 AND Y = 109 else
"110111011111" when X = 28 AND Y = 109 else
"110111011111" when X = 29 AND Y = 109 else
"110111011111" when X = 30 AND Y = 109 else
"110111011111" when X = 31 AND Y = 109 else
"110111011111" when X = 32 AND Y = 109 else
"110111011111" when X = 33 AND Y = 109 else
"110111011111" when X = 34 AND Y = 109 else
"110111011111" when X = 35 AND Y = 109 else
"110111011111" when X = 36 AND Y = 109 else
"110111011111" when X = 37 AND Y = 109 else
"110111011111" when X = 38 AND Y = 109 else
"110111011111" when X = 39 AND Y = 109 else
"110111011111" when X = 40 AND Y = 109 else
"110111011111" when X = 41 AND Y = 109 else
"110111011111" when X = 42 AND Y = 109 else
"110111011111" when X = 43 AND Y = 109 else
"110111011111" when X = 44 AND Y = 109 else
"110111011111" when X = 45 AND Y = 109 else
"110111011111" when X = 46 AND Y = 109 else
"110111011111" when X = 47 AND Y = 109 else
"110111011111" when X = 48 AND Y = 109 else
"110111011111" when X = 49 AND Y = 109 else
"110111011111" when X = 50 AND Y = 109 else
"110111011111" when X = 51 AND Y = 109 else
"110111011111" when X = 52 AND Y = 109 else
"110111011111" when X = 53 AND Y = 109 else
"110111011111" when X = 54 AND Y = 109 else
"110111011111" when X = 55 AND Y = 109 else
"110111011111" when X = 56 AND Y = 109 else
"110111011111" when X = 57 AND Y = 109 else
"110111011111" when X = 58 AND Y = 109 else
"110111011111" when X = 59 AND Y = 109 else
"110111011111" when X = 60 AND Y = 109 else
"110111011111" when X = 61 AND Y = 109 else
"110111011111" when X = 62 AND Y = 109 else
"110111011111" when X = 63 AND Y = 109 else
"110111011111" when X = 64 AND Y = 109 else
"110111011111" when X = 65 AND Y = 109 else
"110111011111" when X = 66 AND Y = 109 else
"110111011111" when X = 67 AND Y = 109 else
"110111011111" when X = 68 AND Y = 109 else
"110111011111" when X = 69 AND Y = 109 else
"111111111111" when X = 70 AND Y = 109 else
"111111111111" when X = 71 AND Y = 109 else
"111111111111" when X = 72 AND Y = 109 else
"111111111111" when X = 73 AND Y = 109 else
"111111111111" when X = 74 AND Y = 109 else
"111111111111" when X = 75 AND Y = 109 else
"111111111111" when X = 76 AND Y = 109 else
"111111111111" when X = 77 AND Y = 109 else
"111111111111" when X = 78 AND Y = 109 else
"111111111111" when X = 79 AND Y = 109 else
"111111111111" when X = 80 AND Y = 109 else
"111111111111" when X = 81 AND Y = 109 else
"111111111111" when X = 82 AND Y = 109 else
"111111111111" when X = 83 AND Y = 109 else
"111111111111" when X = 84 AND Y = 109 else
"111111111111" when X = 85 AND Y = 109 else
"111111111111" when X = 86 AND Y = 109 else
"111111111111" when X = 87 AND Y = 109 else
"111111111111" when X = 88 AND Y = 109 else
"111111111111" when X = 89 AND Y = 109 else
"111111111111" when X = 90 AND Y = 109 else
"111111111111" when X = 91 AND Y = 109 else
"111111111111" when X = 92 AND Y = 109 else
"111111111111" when X = 93 AND Y = 109 else
"111111111111" when X = 94 AND Y = 109 else
"111111111111" when X = 95 AND Y = 109 else
"111111111111" when X = 96 AND Y = 109 else
"111111111111" when X = 97 AND Y = 109 else
"111111111111" when X = 98 AND Y = 109 else
"111111111111" when X = 99 AND Y = 109 else
"111111111111" when X = 100 AND Y = 109 else
"111111111111" when X = 101 AND Y = 109 else
"111111111111" when X = 102 AND Y = 109 else
"111111111111" when X = 103 AND Y = 109 else
"111111111111" when X = 104 AND Y = 109 else
"111111111111" when X = 105 AND Y = 109 else
"111111111111" when X = 106 AND Y = 109 else
"111111111111" when X = 107 AND Y = 109 else
"111111111111" when X = 108 AND Y = 109 else
"111111111111" when X = 109 AND Y = 109 else
"111111111111" when X = 110 AND Y = 109 else
"111111111111" when X = 111 AND Y = 109 else
"111111111111" when X = 112 AND Y = 109 else
"111111111111" when X = 113 AND Y = 109 else
"111111111111" when X = 114 AND Y = 109 else
"111111111111" when X = 115 AND Y = 109 else
"111111111111" when X = 116 AND Y = 109 else
"111111111111" when X = 117 AND Y = 109 else
"111111111111" when X = 118 AND Y = 109 else
"111111111111" when X = 119 AND Y = 109 else
"111111111111" when X = 120 AND Y = 109 else
"111111111111" when X = 121 AND Y = 109 else
"111111111111" when X = 122 AND Y = 109 else
"111111111111" when X = 123 AND Y = 109 else
"111111111111" when X = 124 AND Y = 109 else
"111111111111" when X = 125 AND Y = 109 else
"111111111111" when X = 126 AND Y = 109 else
"111111111111" when X = 127 AND Y = 109 else
"111111111111" when X = 128 AND Y = 109 else
"111111111111" when X = 129 AND Y = 109 else
"111111111111" when X = 130 AND Y = 109 else
"111111111111" when X = 131 AND Y = 109 else
"111111111111" when X = 132 AND Y = 109 else
"111111111111" when X = 133 AND Y = 109 else
"111111111111" when X = 134 AND Y = 109 else
"111111111111" when X = 135 AND Y = 109 else
"111111111111" when X = 136 AND Y = 109 else
"111111111111" when X = 137 AND Y = 109 else
"111111111111" when X = 138 AND Y = 109 else
"111111111111" when X = 139 AND Y = 109 else
"111111111111" when X = 140 AND Y = 109 else
"111111111111" when X = 141 AND Y = 109 else
"111111111111" when X = 142 AND Y = 109 else
"111111111111" when X = 143 AND Y = 109 else
"111111111111" when X = 144 AND Y = 109 else
"111111111111" when X = 145 AND Y = 109 else
"111111111111" when X = 146 AND Y = 109 else
"111111111111" when X = 147 AND Y = 109 else
"111111111111" when X = 148 AND Y = 109 else
"111111111111" when X = 149 AND Y = 109 else
"111111111111" when X = 150 AND Y = 109 else
"111111111111" when X = 151 AND Y = 109 else
"111111111111" when X = 152 AND Y = 109 else
"111111111111" when X = 153 AND Y = 109 else
"111111111111" when X = 154 AND Y = 109 else
"111111111111" when X = 155 AND Y = 109 else
"111111111111" when X = 156 AND Y = 109 else
"111111111111" when X = 157 AND Y = 109 else
"111111111111" when X = 158 AND Y = 109 else
"111111111111" when X = 159 AND Y = 109 else
"110111011111" when X = 160 AND Y = 109 else
"110111011111" when X = 161 AND Y = 109 else
"110111011111" when X = 162 AND Y = 109 else
"110111011111" when X = 163 AND Y = 109 else
"110111011111" when X = 164 AND Y = 109 else
"110111011111" when X = 165 AND Y = 109 else
"110111011111" when X = 166 AND Y = 109 else
"110111011111" when X = 167 AND Y = 109 else
"110111011111" when X = 168 AND Y = 109 else
"110111011111" when X = 169 AND Y = 109 else
"110111011111" when X = 170 AND Y = 109 else
"110111011111" when X = 171 AND Y = 109 else
"110111011111" when X = 172 AND Y = 109 else
"110111011111" when X = 173 AND Y = 109 else
"110111011111" when X = 174 AND Y = 109 else
"110111011111" when X = 175 AND Y = 109 else
"110111011111" when X = 176 AND Y = 109 else
"110111011111" when X = 177 AND Y = 109 else
"110111011111" when X = 178 AND Y = 109 else
"110111011111" when X = 179 AND Y = 109 else
"110111011111" when X = 180 AND Y = 109 else
"110111011111" when X = 181 AND Y = 109 else
"110111011111" when X = 182 AND Y = 109 else
"110111011111" when X = 183 AND Y = 109 else
"110111011111" when X = 184 AND Y = 109 else
"110111011111" when X = 185 AND Y = 109 else
"110111011111" when X = 186 AND Y = 109 else
"110111011111" when X = 187 AND Y = 109 else
"110111011111" when X = 188 AND Y = 109 else
"110111011111" when X = 189 AND Y = 109 else
"110111011111" when X = 190 AND Y = 109 else
"110111011111" when X = 191 AND Y = 109 else
"110111011111" when X = 192 AND Y = 109 else
"110111011111" when X = 193 AND Y = 109 else
"110111011111" when X = 194 AND Y = 109 else
"110111011111" when X = 195 AND Y = 109 else
"110111011111" when X = 196 AND Y = 109 else
"110111011111" when X = 197 AND Y = 109 else
"110111011111" when X = 198 AND Y = 109 else
"110111011111" when X = 199 AND Y = 109 else
"110111011111" when X = 200 AND Y = 109 else
"110111011111" when X = 201 AND Y = 109 else
"110111011111" when X = 202 AND Y = 109 else
"110111011111" when X = 203 AND Y = 109 else
"110111011111" when X = 204 AND Y = 109 else
"111111111111" when X = 205 AND Y = 109 else
"111111111111" when X = 206 AND Y = 109 else
"111111111111" when X = 207 AND Y = 109 else
"111111111111" when X = 208 AND Y = 109 else
"111111111111" when X = 209 AND Y = 109 else
"111111111111" when X = 210 AND Y = 109 else
"111111111111" when X = 211 AND Y = 109 else
"111111111111" when X = 212 AND Y = 109 else
"111111111111" when X = 213 AND Y = 109 else
"111111111111" when X = 214 AND Y = 109 else
"110111011111" when X = 215 AND Y = 109 else
"110111011111" when X = 216 AND Y = 109 else
"110111011111" when X = 217 AND Y = 109 else
"110111011111" when X = 218 AND Y = 109 else
"110111011111" when X = 219 AND Y = 109 else
"110111011111" when X = 220 AND Y = 109 else
"110111011111" when X = 221 AND Y = 109 else
"110111011111" when X = 222 AND Y = 109 else
"110111011111" when X = 223 AND Y = 109 else
"110111011111" when X = 224 AND Y = 109 else
"110111011111" when X = 225 AND Y = 109 else
"110111011111" when X = 226 AND Y = 109 else
"110111011111" when X = 227 AND Y = 109 else
"110111011111" when X = 228 AND Y = 109 else
"110111011111" when X = 229 AND Y = 109 else
"110111011111" when X = 230 AND Y = 109 else
"110111011111" when X = 231 AND Y = 109 else
"110111011111" when X = 232 AND Y = 109 else
"110111011111" when X = 233 AND Y = 109 else
"110111011111" when X = 234 AND Y = 109 else
"110111011111" when X = 235 AND Y = 109 else
"110111011111" when X = 236 AND Y = 109 else
"110111011111" when X = 237 AND Y = 109 else
"110111011111" when X = 238 AND Y = 109 else
"110111011111" when X = 239 AND Y = 109 else
"110111011111" when X = 240 AND Y = 109 else
"110111011111" when X = 241 AND Y = 109 else
"110111011111" when X = 242 AND Y = 109 else
"110111011111" when X = 243 AND Y = 109 else
"110111011111" when X = 244 AND Y = 109 else
"110111011111" when X = 245 AND Y = 109 else
"110111011111" when X = 246 AND Y = 109 else
"110111011111" when X = 247 AND Y = 109 else
"110111011111" when X = 248 AND Y = 109 else
"110111011111" when X = 249 AND Y = 109 else
"110111011111" when X = 250 AND Y = 109 else
"110111011111" when X = 251 AND Y = 109 else
"110111011111" when X = 252 AND Y = 109 else
"110111011111" when X = 253 AND Y = 109 else
"110111011111" when X = 254 AND Y = 109 else
"110111011111" when X = 255 AND Y = 109 else
"110111011111" when X = 256 AND Y = 109 else
"110111011111" when X = 257 AND Y = 109 else
"110111011111" when X = 258 AND Y = 109 else
"110111011111" when X = 259 AND Y = 109 else
"110111011111" when X = 260 AND Y = 109 else
"110111011111" when X = 261 AND Y = 109 else
"110111011111" when X = 262 AND Y = 109 else
"110111011111" when X = 263 AND Y = 109 else
"110111011111" when X = 264 AND Y = 109 else
"110111011111" when X = 265 AND Y = 109 else
"110111011111" when X = 266 AND Y = 109 else
"110111011111" when X = 267 AND Y = 109 else
"110111011111" when X = 268 AND Y = 109 else
"110111011111" when X = 269 AND Y = 109 else
"110111011111" when X = 270 AND Y = 109 else
"110111011111" when X = 271 AND Y = 109 else
"110111011111" when X = 272 AND Y = 109 else
"110111011111" when X = 273 AND Y = 109 else
"110111011111" when X = 274 AND Y = 109 else
"110111011111" when X = 275 AND Y = 109 else
"110111011111" when X = 276 AND Y = 109 else
"110111011111" when X = 277 AND Y = 109 else
"110111011111" when X = 278 AND Y = 109 else
"110111011111" when X = 279 AND Y = 109 else
"111111111111" when X = 280 AND Y = 109 else
"111111111111" when X = 281 AND Y = 109 else
"111111111111" when X = 282 AND Y = 109 else
"111111111111" when X = 283 AND Y = 109 else
"111111111111" when X = 284 AND Y = 109 else
"111111111111" when X = 285 AND Y = 109 else
"111111111111" when X = 286 AND Y = 109 else
"111111111111" when X = 287 AND Y = 109 else
"111111111111" when X = 288 AND Y = 109 else
"111111111111" when X = 289 AND Y = 109 else
"111111111111" when X = 290 AND Y = 109 else
"111111111111" when X = 291 AND Y = 109 else
"111111111111" when X = 292 AND Y = 109 else
"111111111111" when X = 293 AND Y = 109 else
"111111111111" when X = 294 AND Y = 109 else
"111111111111" when X = 295 AND Y = 109 else
"111111111111" when X = 296 AND Y = 109 else
"111111111111" when X = 297 AND Y = 109 else
"111111111111" when X = 298 AND Y = 109 else
"111111111111" when X = 299 AND Y = 109 else
"111111111111" when X = 300 AND Y = 109 else
"111111111111" when X = 301 AND Y = 109 else
"111111111111" when X = 302 AND Y = 109 else
"111111111111" when X = 303 AND Y = 109 else
"111111111111" when X = 304 AND Y = 109 else
"110111011111" when X = 305 AND Y = 109 else
"110111011111" when X = 306 AND Y = 109 else
"110111011111" when X = 307 AND Y = 109 else
"110111011111" when X = 308 AND Y = 109 else
"110111011111" when X = 309 AND Y = 109 else
"110111011111" when X = 310 AND Y = 109 else
"110111011111" when X = 311 AND Y = 109 else
"110111011111" when X = 312 AND Y = 109 else
"110111011111" when X = 313 AND Y = 109 else
"110111011111" when X = 314 AND Y = 109 else
"110111011111" when X = 315 AND Y = 109 else
"110111011111" when X = 316 AND Y = 109 else
"110111011111" when X = 317 AND Y = 109 else
"110111011111" when X = 318 AND Y = 109 else
"110111011111" when X = 319 AND Y = 109 else
"110111011111" when X = 320 AND Y = 109 else
"110111011111" when X = 321 AND Y = 109 else
"110111011111" when X = 322 AND Y = 109 else
"110111011111" when X = 323 AND Y = 109 else
"110111011111" when X = 324 AND Y = 109 else
"100010011101" when X = 0 AND Y = 110 else
"100010011101" when X = 1 AND Y = 110 else
"100010011101" when X = 2 AND Y = 110 else
"100010011101" when X = 3 AND Y = 110 else
"100010011101" when X = 4 AND Y = 110 else
"100010011101" when X = 5 AND Y = 110 else
"100010011101" when X = 6 AND Y = 110 else
"100010011101" when X = 7 AND Y = 110 else
"100010011101" when X = 8 AND Y = 110 else
"100010011101" when X = 9 AND Y = 110 else
"100010011101" when X = 10 AND Y = 110 else
"100010011101" when X = 11 AND Y = 110 else
"100010011101" when X = 12 AND Y = 110 else
"100010011101" when X = 13 AND Y = 110 else
"100010011101" when X = 14 AND Y = 110 else
"100010011101" when X = 15 AND Y = 110 else
"100010011101" when X = 16 AND Y = 110 else
"100010011101" when X = 17 AND Y = 110 else
"100010011101" when X = 18 AND Y = 110 else
"100010011101" when X = 19 AND Y = 110 else
"100010011101" when X = 20 AND Y = 110 else
"100010011101" when X = 21 AND Y = 110 else
"100010011101" when X = 22 AND Y = 110 else
"100010011101" when X = 23 AND Y = 110 else
"100010011101" when X = 24 AND Y = 110 else
"110111011111" when X = 25 AND Y = 110 else
"110111011111" when X = 26 AND Y = 110 else
"110111011111" when X = 27 AND Y = 110 else
"110111011111" when X = 28 AND Y = 110 else
"110111011111" when X = 29 AND Y = 110 else
"110111011111" when X = 30 AND Y = 110 else
"110111011111" when X = 31 AND Y = 110 else
"110111011111" when X = 32 AND Y = 110 else
"110111011111" when X = 33 AND Y = 110 else
"110111011111" when X = 34 AND Y = 110 else
"110111011111" when X = 35 AND Y = 110 else
"110111011111" when X = 36 AND Y = 110 else
"110111011111" when X = 37 AND Y = 110 else
"110111011111" when X = 38 AND Y = 110 else
"110111011111" when X = 39 AND Y = 110 else
"110111011111" when X = 40 AND Y = 110 else
"110111011111" when X = 41 AND Y = 110 else
"110111011111" when X = 42 AND Y = 110 else
"110111011111" when X = 43 AND Y = 110 else
"110111011111" when X = 44 AND Y = 110 else
"110111011111" when X = 45 AND Y = 110 else
"110111011111" when X = 46 AND Y = 110 else
"110111011111" when X = 47 AND Y = 110 else
"110111011111" when X = 48 AND Y = 110 else
"110111011111" when X = 49 AND Y = 110 else
"110111011111" when X = 50 AND Y = 110 else
"110111011111" when X = 51 AND Y = 110 else
"110111011111" when X = 52 AND Y = 110 else
"110111011111" when X = 53 AND Y = 110 else
"110111011111" when X = 54 AND Y = 110 else
"110111011111" when X = 55 AND Y = 110 else
"110111011111" when X = 56 AND Y = 110 else
"110111011111" when X = 57 AND Y = 110 else
"110111011111" when X = 58 AND Y = 110 else
"110111011111" when X = 59 AND Y = 110 else
"110111011111" when X = 60 AND Y = 110 else
"110111011111" when X = 61 AND Y = 110 else
"110111011111" when X = 62 AND Y = 110 else
"110111011111" when X = 63 AND Y = 110 else
"110111011111" when X = 64 AND Y = 110 else
"110111011111" when X = 65 AND Y = 110 else
"110111011111" when X = 66 AND Y = 110 else
"110111011111" when X = 67 AND Y = 110 else
"110111011111" when X = 68 AND Y = 110 else
"110111011111" when X = 69 AND Y = 110 else
"111111111111" when X = 70 AND Y = 110 else
"111111111111" when X = 71 AND Y = 110 else
"111111111111" when X = 72 AND Y = 110 else
"111111111111" when X = 73 AND Y = 110 else
"111111111111" when X = 74 AND Y = 110 else
"111111111111" when X = 75 AND Y = 110 else
"111111111111" when X = 76 AND Y = 110 else
"111111111111" when X = 77 AND Y = 110 else
"111111111111" when X = 78 AND Y = 110 else
"111111111111" when X = 79 AND Y = 110 else
"111111111111" when X = 80 AND Y = 110 else
"111111111111" when X = 81 AND Y = 110 else
"111111111111" when X = 82 AND Y = 110 else
"111111111111" when X = 83 AND Y = 110 else
"111111111111" when X = 84 AND Y = 110 else
"111111111111" when X = 85 AND Y = 110 else
"111111111111" when X = 86 AND Y = 110 else
"111111111111" when X = 87 AND Y = 110 else
"111111111111" when X = 88 AND Y = 110 else
"111111111111" when X = 89 AND Y = 110 else
"111111111111" when X = 90 AND Y = 110 else
"111111111111" when X = 91 AND Y = 110 else
"111111111111" when X = 92 AND Y = 110 else
"111111111111" when X = 93 AND Y = 110 else
"111111111111" when X = 94 AND Y = 110 else
"111111111111" when X = 95 AND Y = 110 else
"111111111111" when X = 96 AND Y = 110 else
"111111111111" when X = 97 AND Y = 110 else
"111111111111" when X = 98 AND Y = 110 else
"111111111111" when X = 99 AND Y = 110 else
"111111111111" when X = 100 AND Y = 110 else
"111111111111" when X = 101 AND Y = 110 else
"111111111111" when X = 102 AND Y = 110 else
"111111111111" when X = 103 AND Y = 110 else
"111111111111" when X = 104 AND Y = 110 else
"111111111111" when X = 105 AND Y = 110 else
"111111111111" when X = 106 AND Y = 110 else
"111111111111" when X = 107 AND Y = 110 else
"111111111111" when X = 108 AND Y = 110 else
"111111111111" when X = 109 AND Y = 110 else
"111111111111" when X = 110 AND Y = 110 else
"111111111111" when X = 111 AND Y = 110 else
"111111111111" when X = 112 AND Y = 110 else
"111111111111" when X = 113 AND Y = 110 else
"111111111111" when X = 114 AND Y = 110 else
"111111111111" when X = 115 AND Y = 110 else
"111111111111" when X = 116 AND Y = 110 else
"111111111111" when X = 117 AND Y = 110 else
"111111111111" when X = 118 AND Y = 110 else
"111111111111" when X = 119 AND Y = 110 else
"111111111111" when X = 120 AND Y = 110 else
"111111111111" when X = 121 AND Y = 110 else
"111111111111" when X = 122 AND Y = 110 else
"111111111111" when X = 123 AND Y = 110 else
"111111111111" when X = 124 AND Y = 110 else
"111111111111" when X = 125 AND Y = 110 else
"111111111111" when X = 126 AND Y = 110 else
"111111111111" when X = 127 AND Y = 110 else
"111111111111" when X = 128 AND Y = 110 else
"111111111111" when X = 129 AND Y = 110 else
"111111111111" when X = 130 AND Y = 110 else
"111111111111" when X = 131 AND Y = 110 else
"111111111111" when X = 132 AND Y = 110 else
"111111111111" when X = 133 AND Y = 110 else
"111111111111" when X = 134 AND Y = 110 else
"111111111111" when X = 135 AND Y = 110 else
"111111111111" when X = 136 AND Y = 110 else
"111111111111" when X = 137 AND Y = 110 else
"111111111111" when X = 138 AND Y = 110 else
"111111111111" when X = 139 AND Y = 110 else
"111111111111" when X = 140 AND Y = 110 else
"111111111111" when X = 141 AND Y = 110 else
"111111111111" when X = 142 AND Y = 110 else
"111111111111" when X = 143 AND Y = 110 else
"111111111111" when X = 144 AND Y = 110 else
"111111111111" when X = 145 AND Y = 110 else
"111111111111" when X = 146 AND Y = 110 else
"111111111111" when X = 147 AND Y = 110 else
"111111111111" when X = 148 AND Y = 110 else
"111111111111" when X = 149 AND Y = 110 else
"111111111111" when X = 150 AND Y = 110 else
"111111111111" when X = 151 AND Y = 110 else
"111111111111" when X = 152 AND Y = 110 else
"111111111111" when X = 153 AND Y = 110 else
"111111111111" when X = 154 AND Y = 110 else
"111111111111" when X = 155 AND Y = 110 else
"111111111111" when X = 156 AND Y = 110 else
"111111111111" when X = 157 AND Y = 110 else
"111111111111" when X = 158 AND Y = 110 else
"111111111111" when X = 159 AND Y = 110 else
"111111111111" when X = 160 AND Y = 110 else
"111111111111" when X = 161 AND Y = 110 else
"111111111111" when X = 162 AND Y = 110 else
"111111111111" when X = 163 AND Y = 110 else
"111111111111" when X = 164 AND Y = 110 else
"111111111111" when X = 165 AND Y = 110 else
"111111111111" when X = 166 AND Y = 110 else
"111111111111" when X = 167 AND Y = 110 else
"111111111111" when X = 168 AND Y = 110 else
"111111111111" when X = 169 AND Y = 110 else
"111111111111" when X = 170 AND Y = 110 else
"111111111111" when X = 171 AND Y = 110 else
"111111111111" when X = 172 AND Y = 110 else
"111111111111" when X = 173 AND Y = 110 else
"111111111111" when X = 174 AND Y = 110 else
"111111111111" when X = 175 AND Y = 110 else
"111111111111" when X = 176 AND Y = 110 else
"111111111111" when X = 177 AND Y = 110 else
"111111111111" when X = 178 AND Y = 110 else
"111111111111" when X = 179 AND Y = 110 else
"111111111111" when X = 180 AND Y = 110 else
"111111111111" when X = 181 AND Y = 110 else
"111111111111" when X = 182 AND Y = 110 else
"111111111111" when X = 183 AND Y = 110 else
"111111111111" when X = 184 AND Y = 110 else
"111111111111" when X = 185 AND Y = 110 else
"111111111111" when X = 186 AND Y = 110 else
"111111111111" when X = 187 AND Y = 110 else
"111111111111" when X = 188 AND Y = 110 else
"111111111111" when X = 189 AND Y = 110 else
"111111111111" when X = 190 AND Y = 110 else
"111111111111" when X = 191 AND Y = 110 else
"111111111111" when X = 192 AND Y = 110 else
"111111111111" when X = 193 AND Y = 110 else
"111111111111" when X = 194 AND Y = 110 else
"111111111111" when X = 195 AND Y = 110 else
"111111111111" when X = 196 AND Y = 110 else
"111111111111" when X = 197 AND Y = 110 else
"111111111111" when X = 198 AND Y = 110 else
"111111111111" when X = 199 AND Y = 110 else
"111111111111" when X = 200 AND Y = 110 else
"111111111111" when X = 201 AND Y = 110 else
"111111111111" when X = 202 AND Y = 110 else
"111111111111" when X = 203 AND Y = 110 else
"111111111111" when X = 204 AND Y = 110 else
"111111111111" when X = 205 AND Y = 110 else
"111111111111" when X = 206 AND Y = 110 else
"111111111111" when X = 207 AND Y = 110 else
"111111111111" when X = 208 AND Y = 110 else
"111111111111" when X = 209 AND Y = 110 else
"110111011111" when X = 210 AND Y = 110 else
"110111011111" when X = 211 AND Y = 110 else
"110111011111" when X = 212 AND Y = 110 else
"110111011111" when X = 213 AND Y = 110 else
"110111011111" when X = 214 AND Y = 110 else
"110111011111" when X = 215 AND Y = 110 else
"110111011111" when X = 216 AND Y = 110 else
"110111011111" when X = 217 AND Y = 110 else
"110111011111" when X = 218 AND Y = 110 else
"110111011111" when X = 219 AND Y = 110 else
"110111011111" when X = 220 AND Y = 110 else
"110111011111" when X = 221 AND Y = 110 else
"110111011111" when X = 222 AND Y = 110 else
"110111011111" when X = 223 AND Y = 110 else
"110111011111" when X = 224 AND Y = 110 else
"110111011111" when X = 225 AND Y = 110 else
"110111011111" when X = 226 AND Y = 110 else
"110111011111" when X = 227 AND Y = 110 else
"110111011111" when X = 228 AND Y = 110 else
"110111011111" when X = 229 AND Y = 110 else
"110111011111" when X = 230 AND Y = 110 else
"110111011111" when X = 231 AND Y = 110 else
"110111011111" when X = 232 AND Y = 110 else
"110111011111" when X = 233 AND Y = 110 else
"110111011111" when X = 234 AND Y = 110 else
"110111011111" when X = 235 AND Y = 110 else
"110111011111" when X = 236 AND Y = 110 else
"110111011111" when X = 237 AND Y = 110 else
"110111011111" when X = 238 AND Y = 110 else
"110111011111" when X = 239 AND Y = 110 else
"110111011111" when X = 240 AND Y = 110 else
"110111011111" when X = 241 AND Y = 110 else
"110111011111" when X = 242 AND Y = 110 else
"110111011111" when X = 243 AND Y = 110 else
"110111011111" when X = 244 AND Y = 110 else
"110111011111" when X = 245 AND Y = 110 else
"110111011111" when X = 246 AND Y = 110 else
"110111011111" when X = 247 AND Y = 110 else
"110111011111" when X = 248 AND Y = 110 else
"110111011111" when X = 249 AND Y = 110 else
"110111011111" when X = 250 AND Y = 110 else
"110111011111" when X = 251 AND Y = 110 else
"110111011111" when X = 252 AND Y = 110 else
"110111011111" when X = 253 AND Y = 110 else
"110111011111" when X = 254 AND Y = 110 else
"110111011111" when X = 255 AND Y = 110 else
"110111011111" when X = 256 AND Y = 110 else
"110111011111" when X = 257 AND Y = 110 else
"110111011111" when X = 258 AND Y = 110 else
"110111011111" when X = 259 AND Y = 110 else
"110111011111" when X = 260 AND Y = 110 else
"110111011111" when X = 261 AND Y = 110 else
"110111011111" when X = 262 AND Y = 110 else
"110111011111" when X = 263 AND Y = 110 else
"110111011111" when X = 264 AND Y = 110 else
"110111011111" when X = 265 AND Y = 110 else
"110111011111" when X = 266 AND Y = 110 else
"110111011111" when X = 267 AND Y = 110 else
"110111011111" when X = 268 AND Y = 110 else
"110111011111" when X = 269 AND Y = 110 else
"110111011111" when X = 270 AND Y = 110 else
"110111011111" when X = 271 AND Y = 110 else
"110111011111" when X = 272 AND Y = 110 else
"110111011111" when X = 273 AND Y = 110 else
"110111011111" when X = 274 AND Y = 110 else
"110111011111" when X = 275 AND Y = 110 else
"110111011111" when X = 276 AND Y = 110 else
"110111011111" when X = 277 AND Y = 110 else
"110111011111" when X = 278 AND Y = 110 else
"110111011111" when X = 279 AND Y = 110 else
"111111111111" when X = 280 AND Y = 110 else
"111111111111" when X = 281 AND Y = 110 else
"111111111111" when X = 282 AND Y = 110 else
"111111111111" when X = 283 AND Y = 110 else
"111111111111" when X = 284 AND Y = 110 else
"111111111111" when X = 285 AND Y = 110 else
"111111111111" when X = 286 AND Y = 110 else
"111111111111" when X = 287 AND Y = 110 else
"111111111111" when X = 288 AND Y = 110 else
"111111111111" when X = 289 AND Y = 110 else
"111111111111" when X = 290 AND Y = 110 else
"111111111111" when X = 291 AND Y = 110 else
"111111111111" when X = 292 AND Y = 110 else
"111111111111" when X = 293 AND Y = 110 else
"111111111111" when X = 294 AND Y = 110 else
"111111111111" when X = 295 AND Y = 110 else
"111111111111" when X = 296 AND Y = 110 else
"111111111111" when X = 297 AND Y = 110 else
"111111111111" when X = 298 AND Y = 110 else
"111111111111" when X = 299 AND Y = 110 else
"111111111111" when X = 300 AND Y = 110 else
"111111111111" when X = 301 AND Y = 110 else
"111111111111" when X = 302 AND Y = 110 else
"111111111111" when X = 303 AND Y = 110 else
"111111111111" when X = 304 AND Y = 110 else
"110111011111" when X = 305 AND Y = 110 else
"110111011111" when X = 306 AND Y = 110 else
"110111011111" when X = 307 AND Y = 110 else
"110111011111" when X = 308 AND Y = 110 else
"110111011111" when X = 309 AND Y = 110 else
"110111011111" when X = 310 AND Y = 110 else
"110111011111" when X = 311 AND Y = 110 else
"110111011111" when X = 312 AND Y = 110 else
"110111011111" when X = 313 AND Y = 110 else
"110111011111" when X = 314 AND Y = 110 else
"110111011111" when X = 315 AND Y = 110 else
"110111011111" when X = 316 AND Y = 110 else
"110111011111" when X = 317 AND Y = 110 else
"110111011111" when X = 318 AND Y = 110 else
"110111011111" when X = 319 AND Y = 110 else
"110111011111" when X = 320 AND Y = 110 else
"110111011111" when X = 321 AND Y = 110 else
"110111011111" when X = 322 AND Y = 110 else
"110111011111" when X = 323 AND Y = 110 else
"110111011111" when X = 324 AND Y = 110 else
"100010011101" when X = 0 AND Y = 111 else
"100010011101" when X = 1 AND Y = 111 else
"100010011101" when X = 2 AND Y = 111 else
"100010011101" when X = 3 AND Y = 111 else
"100010011101" when X = 4 AND Y = 111 else
"100010011101" when X = 5 AND Y = 111 else
"100010011101" when X = 6 AND Y = 111 else
"100010011101" when X = 7 AND Y = 111 else
"100010011101" when X = 8 AND Y = 111 else
"100010011101" when X = 9 AND Y = 111 else
"100010011101" when X = 10 AND Y = 111 else
"100010011101" when X = 11 AND Y = 111 else
"100010011101" when X = 12 AND Y = 111 else
"100010011101" when X = 13 AND Y = 111 else
"100010011101" when X = 14 AND Y = 111 else
"100010011101" when X = 15 AND Y = 111 else
"100010011101" when X = 16 AND Y = 111 else
"100010011101" when X = 17 AND Y = 111 else
"100010011101" when X = 18 AND Y = 111 else
"100010011101" when X = 19 AND Y = 111 else
"100010011101" when X = 20 AND Y = 111 else
"100010011101" when X = 21 AND Y = 111 else
"100010011101" when X = 22 AND Y = 111 else
"100010011101" when X = 23 AND Y = 111 else
"100010011101" when X = 24 AND Y = 111 else
"110111011111" when X = 25 AND Y = 111 else
"110111011111" when X = 26 AND Y = 111 else
"110111011111" when X = 27 AND Y = 111 else
"110111011111" when X = 28 AND Y = 111 else
"110111011111" when X = 29 AND Y = 111 else
"110111011111" when X = 30 AND Y = 111 else
"110111011111" when X = 31 AND Y = 111 else
"110111011111" when X = 32 AND Y = 111 else
"110111011111" when X = 33 AND Y = 111 else
"110111011111" when X = 34 AND Y = 111 else
"110111011111" when X = 35 AND Y = 111 else
"110111011111" when X = 36 AND Y = 111 else
"110111011111" when X = 37 AND Y = 111 else
"110111011111" when X = 38 AND Y = 111 else
"110111011111" when X = 39 AND Y = 111 else
"110111011111" when X = 40 AND Y = 111 else
"110111011111" when X = 41 AND Y = 111 else
"110111011111" when X = 42 AND Y = 111 else
"110111011111" when X = 43 AND Y = 111 else
"110111011111" when X = 44 AND Y = 111 else
"110111011111" when X = 45 AND Y = 111 else
"110111011111" when X = 46 AND Y = 111 else
"110111011111" when X = 47 AND Y = 111 else
"110111011111" when X = 48 AND Y = 111 else
"110111011111" when X = 49 AND Y = 111 else
"110111011111" when X = 50 AND Y = 111 else
"110111011111" when X = 51 AND Y = 111 else
"110111011111" when X = 52 AND Y = 111 else
"110111011111" when X = 53 AND Y = 111 else
"110111011111" when X = 54 AND Y = 111 else
"110111011111" when X = 55 AND Y = 111 else
"110111011111" when X = 56 AND Y = 111 else
"110111011111" when X = 57 AND Y = 111 else
"110111011111" when X = 58 AND Y = 111 else
"110111011111" when X = 59 AND Y = 111 else
"110111011111" when X = 60 AND Y = 111 else
"110111011111" when X = 61 AND Y = 111 else
"110111011111" when X = 62 AND Y = 111 else
"110111011111" when X = 63 AND Y = 111 else
"110111011111" when X = 64 AND Y = 111 else
"110111011111" when X = 65 AND Y = 111 else
"110111011111" when X = 66 AND Y = 111 else
"110111011111" when X = 67 AND Y = 111 else
"110111011111" when X = 68 AND Y = 111 else
"110111011111" when X = 69 AND Y = 111 else
"111111111111" when X = 70 AND Y = 111 else
"111111111111" when X = 71 AND Y = 111 else
"111111111111" when X = 72 AND Y = 111 else
"111111111111" when X = 73 AND Y = 111 else
"111111111111" when X = 74 AND Y = 111 else
"111111111111" when X = 75 AND Y = 111 else
"111111111111" when X = 76 AND Y = 111 else
"111111111111" when X = 77 AND Y = 111 else
"111111111111" when X = 78 AND Y = 111 else
"111111111111" when X = 79 AND Y = 111 else
"111111111111" when X = 80 AND Y = 111 else
"111111111111" when X = 81 AND Y = 111 else
"111111111111" when X = 82 AND Y = 111 else
"111111111111" when X = 83 AND Y = 111 else
"111111111111" when X = 84 AND Y = 111 else
"111111111111" when X = 85 AND Y = 111 else
"111111111111" when X = 86 AND Y = 111 else
"111111111111" when X = 87 AND Y = 111 else
"111111111111" when X = 88 AND Y = 111 else
"111111111111" when X = 89 AND Y = 111 else
"111111111111" when X = 90 AND Y = 111 else
"111111111111" when X = 91 AND Y = 111 else
"111111111111" when X = 92 AND Y = 111 else
"111111111111" when X = 93 AND Y = 111 else
"111111111111" when X = 94 AND Y = 111 else
"111111111111" when X = 95 AND Y = 111 else
"111111111111" when X = 96 AND Y = 111 else
"111111111111" when X = 97 AND Y = 111 else
"111111111111" when X = 98 AND Y = 111 else
"111111111111" when X = 99 AND Y = 111 else
"111111111111" when X = 100 AND Y = 111 else
"111111111111" when X = 101 AND Y = 111 else
"111111111111" when X = 102 AND Y = 111 else
"111111111111" when X = 103 AND Y = 111 else
"111111111111" when X = 104 AND Y = 111 else
"111111111111" when X = 105 AND Y = 111 else
"111111111111" when X = 106 AND Y = 111 else
"111111111111" when X = 107 AND Y = 111 else
"111111111111" when X = 108 AND Y = 111 else
"111111111111" when X = 109 AND Y = 111 else
"111111111111" when X = 110 AND Y = 111 else
"111111111111" when X = 111 AND Y = 111 else
"111111111111" when X = 112 AND Y = 111 else
"111111111111" when X = 113 AND Y = 111 else
"111111111111" when X = 114 AND Y = 111 else
"111111111111" when X = 115 AND Y = 111 else
"111111111111" when X = 116 AND Y = 111 else
"111111111111" when X = 117 AND Y = 111 else
"111111111111" when X = 118 AND Y = 111 else
"111111111111" when X = 119 AND Y = 111 else
"111111111111" when X = 120 AND Y = 111 else
"111111111111" when X = 121 AND Y = 111 else
"111111111111" when X = 122 AND Y = 111 else
"111111111111" when X = 123 AND Y = 111 else
"111111111111" when X = 124 AND Y = 111 else
"111111111111" when X = 125 AND Y = 111 else
"111111111111" when X = 126 AND Y = 111 else
"111111111111" when X = 127 AND Y = 111 else
"111111111111" when X = 128 AND Y = 111 else
"111111111111" when X = 129 AND Y = 111 else
"111111111111" when X = 130 AND Y = 111 else
"111111111111" when X = 131 AND Y = 111 else
"111111111111" when X = 132 AND Y = 111 else
"111111111111" when X = 133 AND Y = 111 else
"111111111111" when X = 134 AND Y = 111 else
"111111111111" when X = 135 AND Y = 111 else
"111111111111" when X = 136 AND Y = 111 else
"111111111111" when X = 137 AND Y = 111 else
"111111111111" when X = 138 AND Y = 111 else
"111111111111" when X = 139 AND Y = 111 else
"111111111111" when X = 140 AND Y = 111 else
"111111111111" when X = 141 AND Y = 111 else
"111111111111" when X = 142 AND Y = 111 else
"111111111111" when X = 143 AND Y = 111 else
"111111111111" when X = 144 AND Y = 111 else
"111111111111" when X = 145 AND Y = 111 else
"111111111111" when X = 146 AND Y = 111 else
"111111111111" when X = 147 AND Y = 111 else
"111111111111" when X = 148 AND Y = 111 else
"111111111111" when X = 149 AND Y = 111 else
"111111111111" when X = 150 AND Y = 111 else
"111111111111" when X = 151 AND Y = 111 else
"111111111111" when X = 152 AND Y = 111 else
"111111111111" when X = 153 AND Y = 111 else
"111111111111" when X = 154 AND Y = 111 else
"111111111111" when X = 155 AND Y = 111 else
"111111111111" when X = 156 AND Y = 111 else
"111111111111" when X = 157 AND Y = 111 else
"111111111111" when X = 158 AND Y = 111 else
"111111111111" when X = 159 AND Y = 111 else
"111111111111" when X = 160 AND Y = 111 else
"111111111111" when X = 161 AND Y = 111 else
"111111111111" when X = 162 AND Y = 111 else
"111111111111" when X = 163 AND Y = 111 else
"111111111111" when X = 164 AND Y = 111 else
"111111111111" when X = 165 AND Y = 111 else
"111111111111" when X = 166 AND Y = 111 else
"111111111111" when X = 167 AND Y = 111 else
"111111111111" when X = 168 AND Y = 111 else
"111111111111" when X = 169 AND Y = 111 else
"111111111111" when X = 170 AND Y = 111 else
"111111111111" when X = 171 AND Y = 111 else
"111111111111" when X = 172 AND Y = 111 else
"111111111111" when X = 173 AND Y = 111 else
"111111111111" when X = 174 AND Y = 111 else
"111111111111" when X = 175 AND Y = 111 else
"111111111111" when X = 176 AND Y = 111 else
"111111111111" when X = 177 AND Y = 111 else
"111111111111" when X = 178 AND Y = 111 else
"111111111111" when X = 179 AND Y = 111 else
"111111111111" when X = 180 AND Y = 111 else
"111111111111" when X = 181 AND Y = 111 else
"111111111111" when X = 182 AND Y = 111 else
"111111111111" when X = 183 AND Y = 111 else
"111111111111" when X = 184 AND Y = 111 else
"111111111111" when X = 185 AND Y = 111 else
"111111111111" when X = 186 AND Y = 111 else
"111111111111" when X = 187 AND Y = 111 else
"111111111111" when X = 188 AND Y = 111 else
"111111111111" when X = 189 AND Y = 111 else
"111111111111" when X = 190 AND Y = 111 else
"111111111111" when X = 191 AND Y = 111 else
"111111111111" when X = 192 AND Y = 111 else
"111111111111" when X = 193 AND Y = 111 else
"111111111111" when X = 194 AND Y = 111 else
"111111111111" when X = 195 AND Y = 111 else
"111111111111" when X = 196 AND Y = 111 else
"111111111111" when X = 197 AND Y = 111 else
"111111111111" when X = 198 AND Y = 111 else
"111111111111" when X = 199 AND Y = 111 else
"111111111111" when X = 200 AND Y = 111 else
"111111111111" when X = 201 AND Y = 111 else
"111111111111" when X = 202 AND Y = 111 else
"111111111111" when X = 203 AND Y = 111 else
"111111111111" when X = 204 AND Y = 111 else
"111111111111" when X = 205 AND Y = 111 else
"111111111111" when X = 206 AND Y = 111 else
"111111111111" when X = 207 AND Y = 111 else
"111111111111" when X = 208 AND Y = 111 else
"111111111111" when X = 209 AND Y = 111 else
"110111011111" when X = 210 AND Y = 111 else
"110111011111" when X = 211 AND Y = 111 else
"110111011111" when X = 212 AND Y = 111 else
"110111011111" when X = 213 AND Y = 111 else
"110111011111" when X = 214 AND Y = 111 else
"110111011111" when X = 215 AND Y = 111 else
"110111011111" when X = 216 AND Y = 111 else
"110111011111" when X = 217 AND Y = 111 else
"110111011111" when X = 218 AND Y = 111 else
"110111011111" when X = 219 AND Y = 111 else
"110111011111" when X = 220 AND Y = 111 else
"110111011111" when X = 221 AND Y = 111 else
"110111011111" when X = 222 AND Y = 111 else
"110111011111" when X = 223 AND Y = 111 else
"110111011111" when X = 224 AND Y = 111 else
"110111011111" when X = 225 AND Y = 111 else
"110111011111" when X = 226 AND Y = 111 else
"110111011111" when X = 227 AND Y = 111 else
"110111011111" when X = 228 AND Y = 111 else
"110111011111" when X = 229 AND Y = 111 else
"110111011111" when X = 230 AND Y = 111 else
"110111011111" when X = 231 AND Y = 111 else
"110111011111" when X = 232 AND Y = 111 else
"110111011111" when X = 233 AND Y = 111 else
"110111011111" when X = 234 AND Y = 111 else
"110111011111" when X = 235 AND Y = 111 else
"110111011111" when X = 236 AND Y = 111 else
"110111011111" when X = 237 AND Y = 111 else
"110111011111" when X = 238 AND Y = 111 else
"110111011111" when X = 239 AND Y = 111 else
"110111011111" when X = 240 AND Y = 111 else
"110111011111" when X = 241 AND Y = 111 else
"110111011111" when X = 242 AND Y = 111 else
"110111011111" when X = 243 AND Y = 111 else
"110111011111" when X = 244 AND Y = 111 else
"110111011111" when X = 245 AND Y = 111 else
"110111011111" when X = 246 AND Y = 111 else
"110111011111" when X = 247 AND Y = 111 else
"110111011111" when X = 248 AND Y = 111 else
"110111011111" when X = 249 AND Y = 111 else
"110111011111" when X = 250 AND Y = 111 else
"110111011111" when X = 251 AND Y = 111 else
"110111011111" when X = 252 AND Y = 111 else
"110111011111" when X = 253 AND Y = 111 else
"110111011111" when X = 254 AND Y = 111 else
"110111011111" when X = 255 AND Y = 111 else
"110111011111" when X = 256 AND Y = 111 else
"110111011111" when X = 257 AND Y = 111 else
"110111011111" when X = 258 AND Y = 111 else
"110111011111" when X = 259 AND Y = 111 else
"110111011111" when X = 260 AND Y = 111 else
"110111011111" when X = 261 AND Y = 111 else
"110111011111" when X = 262 AND Y = 111 else
"110111011111" when X = 263 AND Y = 111 else
"110111011111" when X = 264 AND Y = 111 else
"110111011111" when X = 265 AND Y = 111 else
"110111011111" when X = 266 AND Y = 111 else
"110111011111" when X = 267 AND Y = 111 else
"110111011111" when X = 268 AND Y = 111 else
"110111011111" when X = 269 AND Y = 111 else
"110111011111" when X = 270 AND Y = 111 else
"110111011111" when X = 271 AND Y = 111 else
"110111011111" when X = 272 AND Y = 111 else
"110111011111" when X = 273 AND Y = 111 else
"110111011111" when X = 274 AND Y = 111 else
"110111011111" when X = 275 AND Y = 111 else
"110111011111" when X = 276 AND Y = 111 else
"110111011111" when X = 277 AND Y = 111 else
"110111011111" when X = 278 AND Y = 111 else
"110111011111" when X = 279 AND Y = 111 else
"111111111111" when X = 280 AND Y = 111 else
"111111111111" when X = 281 AND Y = 111 else
"111111111111" when X = 282 AND Y = 111 else
"111111111111" when X = 283 AND Y = 111 else
"111111111111" when X = 284 AND Y = 111 else
"111111111111" when X = 285 AND Y = 111 else
"111111111111" when X = 286 AND Y = 111 else
"111111111111" when X = 287 AND Y = 111 else
"111111111111" when X = 288 AND Y = 111 else
"111111111111" when X = 289 AND Y = 111 else
"111111111111" when X = 290 AND Y = 111 else
"111111111111" when X = 291 AND Y = 111 else
"111111111111" when X = 292 AND Y = 111 else
"111111111111" when X = 293 AND Y = 111 else
"111111111111" when X = 294 AND Y = 111 else
"111111111111" when X = 295 AND Y = 111 else
"111111111111" when X = 296 AND Y = 111 else
"111111111111" when X = 297 AND Y = 111 else
"111111111111" when X = 298 AND Y = 111 else
"111111111111" when X = 299 AND Y = 111 else
"111111111111" when X = 300 AND Y = 111 else
"111111111111" when X = 301 AND Y = 111 else
"111111111111" when X = 302 AND Y = 111 else
"111111111111" when X = 303 AND Y = 111 else
"111111111111" when X = 304 AND Y = 111 else
"110111011111" when X = 305 AND Y = 111 else
"110111011111" when X = 306 AND Y = 111 else
"110111011111" when X = 307 AND Y = 111 else
"110111011111" when X = 308 AND Y = 111 else
"110111011111" when X = 309 AND Y = 111 else
"110111011111" when X = 310 AND Y = 111 else
"110111011111" when X = 311 AND Y = 111 else
"110111011111" when X = 312 AND Y = 111 else
"110111011111" when X = 313 AND Y = 111 else
"110111011111" when X = 314 AND Y = 111 else
"110111011111" when X = 315 AND Y = 111 else
"110111011111" when X = 316 AND Y = 111 else
"110111011111" when X = 317 AND Y = 111 else
"110111011111" when X = 318 AND Y = 111 else
"110111011111" when X = 319 AND Y = 111 else
"110111011111" when X = 320 AND Y = 111 else
"110111011111" when X = 321 AND Y = 111 else
"110111011111" when X = 322 AND Y = 111 else
"110111011111" when X = 323 AND Y = 111 else
"110111011111" when X = 324 AND Y = 111 else
"100010011101" when X = 0 AND Y = 112 else
"100010011101" when X = 1 AND Y = 112 else
"100010011101" when X = 2 AND Y = 112 else
"100010011101" when X = 3 AND Y = 112 else
"100010011101" when X = 4 AND Y = 112 else
"100010011101" when X = 5 AND Y = 112 else
"100010011101" when X = 6 AND Y = 112 else
"100010011101" when X = 7 AND Y = 112 else
"100010011101" when X = 8 AND Y = 112 else
"100010011101" when X = 9 AND Y = 112 else
"100010011101" when X = 10 AND Y = 112 else
"100010011101" when X = 11 AND Y = 112 else
"100010011101" when X = 12 AND Y = 112 else
"100010011101" when X = 13 AND Y = 112 else
"100010011101" when X = 14 AND Y = 112 else
"100010011101" when X = 15 AND Y = 112 else
"100010011101" when X = 16 AND Y = 112 else
"100010011101" when X = 17 AND Y = 112 else
"100010011101" when X = 18 AND Y = 112 else
"100010011101" when X = 19 AND Y = 112 else
"100010011101" when X = 20 AND Y = 112 else
"100010011101" when X = 21 AND Y = 112 else
"100010011101" when X = 22 AND Y = 112 else
"100010011101" when X = 23 AND Y = 112 else
"100010011101" when X = 24 AND Y = 112 else
"110111011111" when X = 25 AND Y = 112 else
"110111011111" when X = 26 AND Y = 112 else
"110111011111" when X = 27 AND Y = 112 else
"110111011111" when X = 28 AND Y = 112 else
"110111011111" when X = 29 AND Y = 112 else
"110111011111" when X = 30 AND Y = 112 else
"110111011111" when X = 31 AND Y = 112 else
"110111011111" when X = 32 AND Y = 112 else
"110111011111" when X = 33 AND Y = 112 else
"110111011111" when X = 34 AND Y = 112 else
"110111011111" when X = 35 AND Y = 112 else
"110111011111" when X = 36 AND Y = 112 else
"110111011111" when X = 37 AND Y = 112 else
"110111011111" when X = 38 AND Y = 112 else
"110111011111" when X = 39 AND Y = 112 else
"110111011111" when X = 40 AND Y = 112 else
"110111011111" when X = 41 AND Y = 112 else
"110111011111" when X = 42 AND Y = 112 else
"110111011111" when X = 43 AND Y = 112 else
"110111011111" when X = 44 AND Y = 112 else
"110111011111" when X = 45 AND Y = 112 else
"110111011111" when X = 46 AND Y = 112 else
"110111011111" when X = 47 AND Y = 112 else
"110111011111" when X = 48 AND Y = 112 else
"110111011111" when X = 49 AND Y = 112 else
"110111011111" when X = 50 AND Y = 112 else
"110111011111" when X = 51 AND Y = 112 else
"110111011111" when X = 52 AND Y = 112 else
"110111011111" when X = 53 AND Y = 112 else
"110111011111" when X = 54 AND Y = 112 else
"110111011111" when X = 55 AND Y = 112 else
"110111011111" when X = 56 AND Y = 112 else
"110111011111" when X = 57 AND Y = 112 else
"110111011111" when X = 58 AND Y = 112 else
"110111011111" when X = 59 AND Y = 112 else
"110111011111" when X = 60 AND Y = 112 else
"110111011111" when X = 61 AND Y = 112 else
"110111011111" when X = 62 AND Y = 112 else
"110111011111" when X = 63 AND Y = 112 else
"110111011111" when X = 64 AND Y = 112 else
"110111011111" when X = 65 AND Y = 112 else
"110111011111" when X = 66 AND Y = 112 else
"110111011111" when X = 67 AND Y = 112 else
"110111011111" when X = 68 AND Y = 112 else
"110111011111" when X = 69 AND Y = 112 else
"111111111111" when X = 70 AND Y = 112 else
"111111111111" when X = 71 AND Y = 112 else
"111111111111" when X = 72 AND Y = 112 else
"111111111111" when X = 73 AND Y = 112 else
"111111111111" when X = 74 AND Y = 112 else
"111111111111" when X = 75 AND Y = 112 else
"111111111111" when X = 76 AND Y = 112 else
"111111111111" when X = 77 AND Y = 112 else
"111111111111" when X = 78 AND Y = 112 else
"111111111111" when X = 79 AND Y = 112 else
"111111111111" when X = 80 AND Y = 112 else
"111111111111" when X = 81 AND Y = 112 else
"111111111111" when X = 82 AND Y = 112 else
"111111111111" when X = 83 AND Y = 112 else
"111111111111" when X = 84 AND Y = 112 else
"111111111111" when X = 85 AND Y = 112 else
"111111111111" when X = 86 AND Y = 112 else
"111111111111" when X = 87 AND Y = 112 else
"111111111111" when X = 88 AND Y = 112 else
"111111111111" when X = 89 AND Y = 112 else
"111111111111" when X = 90 AND Y = 112 else
"111111111111" when X = 91 AND Y = 112 else
"111111111111" when X = 92 AND Y = 112 else
"111111111111" when X = 93 AND Y = 112 else
"111111111111" when X = 94 AND Y = 112 else
"111111111111" when X = 95 AND Y = 112 else
"111111111111" when X = 96 AND Y = 112 else
"111111111111" when X = 97 AND Y = 112 else
"111111111111" when X = 98 AND Y = 112 else
"111111111111" when X = 99 AND Y = 112 else
"111111111111" when X = 100 AND Y = 112 else
"111111111111" when X = 101 AND Y = 112 else
"111111111111" when X = 102 AND Y = 112 else
"111111111111" when X = 103 AND Y = 112 else
"111111111111" when X = 104 AND Y = 112 else
"111111111111" when X = 105 AND Y = 112 else
"111111111111" when X = 106 AND Y = 112 else
"111111111111" when X = 107 AND Y = 112 else
"111111111111" when X = 108 AND Y = 112 else
"111111111111" when X = 109 AND Y = 112 else
"111111111111" when X = 110 AND Y = 112 else
"111111111111" when X = 111 AND Y = 112 else
"111111111111" when X = 112 AND Y = 112 else
"111111111111" when X = 113 AND Y = 112 else
"111111111111" when X = 114 AND Y = 112 else
"111111111111" when X = 115 AND Y = 112 else
"111111111111" when X = 116 AND Y = 112 else
"111111111111" when X = 117 AND Y = 112 else
"111111111111" when X = 118 AND Y = 112 else
"111111111111" when X = 119 AND Y = 112 else
"111111111111" when X = 120 AND Y = 112 else
"111111111111" when X = 121 AND Y = 112 else
"111111111111" when X = 122 AND Y = 112 else
"111111111111" when X = 123 AND Y = 112 else
"111111111111" when X = 124 AND Y = 112 else
"111111111111" when X = 125 AND Y = 112 else
"111111111111" when X = 126 AND Y = 112 else
"111111111111" when X = 127 AND Y = 112 else
"111111111111" when X = 128 AND Y = 112 else
"111111111111" when X = 129 AND Y = 112 else
"111111111111" when X = 130 AND Y = 112 else
"111111111111" when X = 131 AND Y = 112 else
"111111111111" when X = 132 AND Y = 112 else
"111111111111" when X = 133 AND Y = 112 else
"111111111111" when X = 134 AND Y = 112 else
"111111111111" when X = 135 AND Y = 112 else
"111111111111" when X = 136 AND Y = 112 else
"111111111111" when X = 137 AND Y = 112 else
"111111111111" when X = 138 AND Y = 112 else
"111111111111" when X = 139 AND Y = 112 else
"111111111111" when X = 140 AND Y = 112 else
"111111111111" when X = 141 AND Y = 112 else
"111111111111" when X = 142 AND Y = 112 else
"111111111111" when X = 143 AND Y = 112 else
"111111111111" when X = 144 AND Y = 112 else
"111111111111" when X = 145 AND Y = 112 else
"111111111111" when X = 146 AND Y = 112 else
"111111111111" when X = 147 AND Y = 112 else
"111111111111" when X = 148 AND Y = 112 else
"111111111111" when X = 149 AND Y = 112 else
"111111111111" when X = 150 AND Y = 112 else
"111111111111" when X = 151 AND Y = 112 else
"111111111111" when X = 152 AND Y = 112 else
"111111111111" when X = 153 AND Y = 112 else
"111111111111" when X = 154 AND Y = 112 else
"111111111111" when X = 155 AND Y = 112 else
"111111111111" when X = 156 AND Y = 112 else
"111111111111" when X = 157 AND Y = 112 else
"111111111111" when X = 158 AND Y = 112 else
"111111111111" when X = 159 AND Y = 112 else
"111111111111" when X = 160 AND Y = 112 else
"111111111111" when X = 161 AND Y = 112 else
"111111111111" when X = 162 AND Y = 112 else
"111111111111" when X = 163 AND Y = 112 else
"111111111111" when X = 164 AND Y = 112 else
"111111111111" when X = 165 AND Y = 112 else
"111111111111" when X = 166 AND Y = 112 else
"111111111111" when X = 167 AND Y = 112 else
"111111111111" when X = 168 AND Y = 112 else
"111111111111" when X = 169 AND Y = 112 else
"111111111111" when X = 170 AND Y = 112 else
"111111111111" when X = 171 AND Y = 112 else
"111111111111" when X = 172 AND Y = 112 else
"111111111111" when X = 173 AND Y = 112 else
"111111111111" when X = 174 AND Y = 112 else
"111111111111" when X = 175 AND Y = 112 else
"111111111111" when X = 176 AND Y = 112 else
"111111111111" when X = 177 AND Y = 112 else
"111111111111" when X = 178 AND Y = 112 else
"111111111111" when X = 179 AND Y = 112 else
"111111111111" when X = 180 AND Y = 112 else
"111111111111" when X = 181 AND Y = 112 else
"111111111111" when X = 182 AND Y = 112 else
"111111111111" when X = 183 AND Y = 112 else
"111111111111" when X = 184 AND Y = 112 else
"111111111111" when X = 185 AND Y = 112 else
"111111111111" when X = 186 AND Y = 112 else
"111111111111" when X = 187 AND Y = 112 else
"111111111111" when X = 188 AND Y = 112 else
"111111111111" when X = 189 AND Y = 112 else
"111111111111" when X = 190 AND Y = 112 else
"111111111111" when X = 191 AND Y = 112 else
"111111111111" when X = 192 AND Y = 112 else
"111111111111" when X = 193 AND Y = 112 else
"111111111111" when X = 194 AND Y = 112 else
"111111111111" when X = 195 AND Y = 112 else
"111111111111" when X = 196 AND Y = 112 else
"111111111111" when X = 197 AND Y = 112 else
"111111111111" when X = 198 AND Y = 112 else
"111111111111" when X = 199 AND Y = 112 else
"111111111111" when X = 200 AND Y = 112 else
"111111111111" when X = 201 AND Y = 112 else
"111111111111" when X = 202 AND Y = 112 else
"111111111111" when X = 203 AND Y = 112 else
"111111111111" when X = 204 AND Y = 112 else
"111111111111" when X = 205 AND Y = 112 else
"111111111111" when X = 206 AND Y = 112 else
"111111111111" when X = 207 AND Y = 112 else
"111111111111" when X = 208 AND Y = 112 else
"111111111111" when X = 209 AND Y = 112 else
"110111011111" when X = 210 AND Y = 112 else
"110111011111" when X = 211 AND Y = 112 else
"110111011111" when X = 212 AND Y = 112 else
"110111011111" when X = 213 AND Y = 112 else
"110111011111" when X = 214 AND Y = 112 else
"110111011111" when X = 215 AND Y = 112 else
"110111011111" when X = 216 AND Y = 112 else
"110111011111" when X = 217 AND Y = 112 else
"110111011111" when X = 218 AND Y = 112 else
"110111011111" when X = 219 AND Y = 112 else
"110111011111" when X = 220 AND Y = 112 else
"110111011111" when X = 221 AND Y = 112 else
"110111011111" when X = 222 AND Y = 112 else
"110111011111" when X = 223 AND Y = 112 else
"110111011111" when X = 224 AND Y = 112 else
"110111011111" when X = 225 AND Y = 112 else
"110111011111" when X = 226 AND Y = 112 else
"110111011111" when X = 227 AND Y = 112 else
"110111011111" when X = 228 AND Y = 112 else
"110111011111" when X = 229 AND Y = 112 else
"110111011111" when X = 230 AND Y = 112 else
"110111011111" when X = 231 AND Y = 112 else
"110111011111" when X = 232 AND Y = 112 else
"110111011111" when X = 233 AND Y = 112 else
"110111011111" when X = 234 AND Y = 112 else
"110111011111" when X = 235 AND Y = 112 else
"110111011111" when X = 236 AND Y = 112 else
"110111011111" when X = 237 AND Y = 112 else
"110111011111" when X = 238 AND Y = 112 else
"110111011111" when X = 239 AND Y = 112 else
"110111011111" when X = 240 AND Y = 112 else
"110111011111" when X = 241 AND Y = 112 else
"110111011111" when X = 242 AND Y = 112 else
"110111011111" when X = 243 AND Y = 112 else
"110111011111" when X = 244 AND Y = 112 else
"110111011111" when X = 245 AND Y = 112 else
"110111011111" when X = 246 AND Y = 112 else
"110111011111" when X = 247 AND Y = 112 else
"110111011111" when X = 248 AND Y = 112 else
"110111011111" when X = 249 AND Y = 112 else
"110111011111" when X = 250 AND Y = 112 else
"110111011111" when X = 251 AND Y = 112 else
"110111011111" when X = 252 AND Y = 112 else
"110111011111" when X = 253 AND Y = 112 else
"110111011111" when X = 254 AND Y = 112 else
"110111011111" when X = 255 AND Y = 112 else
"110111011111" when X = 256 AND Y = 112 else
"110111011111" when X = 257 AND Y = 112 else
"110111011111" when X = 258 AND Y = 112 else
"110111011111" when X = 259 AND Y = 112 else
"110111011111" when X = 260 AND Y = 112 else
"110111011111" when X = 261 AND Y = 112 else
"110111011111" when X = 262 AND Y = 112 else
"110111011111" when X = 263 AND Y = 112 else
"110111011111" when X = 264 AND Y = 112 else
"110111011111" when X = 265 AND Y = 112 else
"110111011111" when X = 266 AND Y = 112 else
"110111011111" when X = 267 AND Y = 112 else
"110111011111" when X = 268 AND Y = 112 else
"110111011111" when X = 269 AND Y = 112 else
"110111011111" when X = 270 AND Y = 112 else
"110111011111" when X = 271 AND Y = 112 else
"110111011111" when X = 272 AND Y = 112 else
"110111011111" when X = 273 AND Y = 112 else
"110111011111" when X = 274 AND Y = 112 else
"110111011111" when X = 275 AND Y = 112 else
"110111011111" when X = 276 AND Y = 112 else
"110111011111" when X = 277 AND Y = 112 else
"110111011111" when X = 278 AND Y = 112 else
"110111011111" when X = 279 AND Y = 112 else
"111111111111" when X = 280 AND Y = 112 else
"111111111111" when X = 281 AND Y = 112 else
"111111111111" when X = 282 AND Y = 112 else
"111111111111" when X = 283 AND Y = 112 else
"111111111111" when X = 284 AND Y = 112 else
"111111111111" when X = 285 AND Y = 112 else
"111111111111" when X = 286 AND Y = 112 else
"111111111111" when X = 287 AND Y = 112 else
"111111111111" when X = 288 AND Y = 112 else
"111111111111" when X = 289 AND Y = 112 else
"111111111111" when X = 290 AND Y = 112 else
"111111111111" when X = 291 AND Y = 112 else
"111111111111" when X = 292 AND Y = 112 else
"111111111111" when X = 293 AND Y = 112 else
"111111111111" when X = 294 AND Y = 112 else
"111111111111" when X = 295 AND Y = 112 else
"111111111111" when X = 296 AND Y = 112 else
"111111111111" when X = 297 AND Y = 112 else
"111111111111" when X = 298 AND Y = 112 else
"111111111111" when X = 299 AND Y = 112 else
"111111111111" when X = 300 AND Y = 112 else
"111111111111" when X = 301 AND Y = 112 else
"111111111111" when X = 302 AND Y = 112 else
"111111111111" when X = 303 AND Y = 112 else
"111111111111" when X = 304 AND Y = 112 else
"110111011111" when X = 305 AND Y = 112 else
"110111011111" when X = 306 AND Y = 112 else
"110111011111" when X = 307 AND Y = 112 else
"110111011111" when X = 308 AND Y = 112 else
"110111011111" when X = 309 AND Y = 112 else
"110111011111" when X = 310 AND Y = 112 else
"110111011111" when X = 311 AND Y = 112 else
"110111011111" when X = 312 AND Y = 112 else
"110111011111" when X = 313 AND Y = 112 else
"110111011111" when X = 314 AND Y = 112 else
"110111011111" when X = 315 AND Y = 112 else
"110111011111" when X = 316 AND Y = 112 else
"110111011111" when X = 317 AND Y = 112 else
"110111011111" when X = 318 AND Y = 112 else
"110111011111" when X = 319 AND Y = 112 else
"110111011111" when X = 320 AND Y = 112 else
"110111011111" when X = 321 AND Y = 112 else
"110111011111" when X = 322 AND Y = 112 else
"110111011111" when X = 323 AND Y = 112 else
"110111011111" when X = 324 AND Y = 112 else
"100010011101" when X = 0 AND Y = 113 else
"100010011101" when X = 1 AND Y = 113 else
"100010011101" when X = 2 AND Y = 113 else
"100010011101" when X = 3 AND Y = 113 else
"100010011101" when X = 4 AND Y = 113 else
"100010011101" when X = 5 AND Y = 113 else
"100010011101" when X = 6 AND Y = 113 else
"100010011101" when X = 7 AND Y = 113 else
"100010011101" when X = 8 AND Y = 113 else
"100010011101" when X = 9 AND Y = 113 else
"100010011101" when X = 10 AND Y = 113 else
"100010011101" when X = 11 AND Y = 113 else
"100010011101" when X = 12 AND Y = 113 else
"100010011101" when X = 13 AND Y = 113 else
"100010011101" when X = 14 AND Y = 113 else
"100010011101" when X = 15 AND Y = 113 else
"100010011101" when X = 16 AND Y = 113 else
"100010011101" when X = 17 AND Y = 113 else
"100010011101" when X = 18 AND Y = 113 else
"100010011101" when X = 19 AND Y = 113 else
"100010011101" when X = 20 AND Y = 113 else
"100010011101" when X = 21 AND Y = 113 else
"100010011101" when X = 22 AND Y = 113 else
"100010011101" when X = 23 AND Y = 113 else
"100010011101" when X = 24 AND Y = 113 else
"110111011111" when X = 25 AND Y = 113 else
"110111011111" when X = 26 AND Y = 113 else
"110111011111" when X = 27 AND Y = 113 else
"110111011111" when X = 28 AND Y = 113 else
"110111011111" when X = 29 AND Y = 113 else
"110111011111" when X = 30 AND Y = 113 else
"110111011111" when X = 31 AND Y = 113 else
"110111011111" when X = 32 AND Y = 113 else
"110111011111" when X = 33 AND Y = 113 else
"110111011111" when X = 34 AND Y = 113 else
"110111011111" when X = 35 AND Y = 113 else
"110111011111" when X = 36 AND Y = 113 else
"110111011111" when X = 37 AND Y = 113 else
"110111011111" when X = 38 AND Y = 113 else
"110111011111" when X = 39 AND Y = 113 else
"110111011111" when X = 40 AND Y = 113 else
"110111011111" when X = 41 AND Y = 113 else
"110111011111" when X = 42 AND Y = 113 else
"110111011111" when X = 43 AND Y = 113 else
"110111011111" when X = 44 AND Y = 113 else
"110111011111" when X = 45 AND Y = 113 else
"110111011111" when X = 46 AND Y = 113 else
"110111011111" when X = 47 AND Y = 113 else
"110111011111" when X = 48 AND Y = 113 else
"110111011111" when X = 49 AND Y = 113 else
"110111011111" when X = 50 AND Y = 113 else
"110111011111" when X = 51 AND Y = 113 else
"110111011111" when X = 52 AND Y = 113 else
"110111011111" when X = 53 AND Y = 113 else
"110111011111" when X = 54 AND Y = 113 else
"110111011111" when X = 55 AND Y = 113 else
"110111011111" when X = 56 AND Y = 113 else
"110111011111" when X = 57 AND Y = 113 else
"110111011111" when X = 58 AND Y = 113 else
"110111011111" when X = 59 AND Y = 113 else
"110111011111" when X = 60 AND Y = 113 else
"110111011111" when X = 61 AND Y = 113 else
"110111011111" when X = 62 AND Y = 113 else
"110111011111" when X = 63 AND Y = 113 else
"110111011111" when X = 64 AND Y = 113 else
"110111011111" when X = 65 AND Y = 113 else
"110111011111" when X = 66 AND Y = 113 else
"110111011111" when X = 67 AND Y = 113 else
"110111011111" when X = 68 AND Y = 113 else
"110111011111" when X = 69 AND Y = 113 else
"111111111111" when X = 70 AND Y = 113 else
"111111111111" when X = 71 AND Y = 113 else
"111111111111" when X = 72 AND Y = 113 else
"111111111111" when X = 73 AND Y = 113 else
"111111111111" when X = 74 AND Y = 113 else
"111111111111" when X = 75 AND Y = 113 else
"111111111111" when X = 76 AND Y = 113 else
"111111111111" when X = 77 AND Y = 113 else
"111111111111" when X = 78 AND Y = 113 else
"111111111111" when X = 79 AND Y = 113 else
"111111111111" when X = 80 AND Y = 113 else
"111111111111" when X = 81 AND Y = 113 else
"111111111111" when X = 82 AND Y = 113 else
"111111111111" when X = 83 AND Y = 113 else
"111111111111" when X = 84 AND Y = 113 else
"111111111111" when X = 85 AND Y = 113 else
"111111111111" when X = 86 AND Y = 113 else
"111111111111" when X = 87 AND Y = 113 else
"111111111111" when X = 88 AND Y = 113 else
"111111111111" when X = 89 AND Y = 113 else
"111111111111" when X = 90 AND Y = 113 else
"111111111111" when X = 91 AND Y = 113 else
"111111111111" when X = 92 AND Y = 113 else
"111111111111" when X = 93 AND Y = 113 else
"111111111111" when X = 94 AND Y = 113 else
"111111111111" when X = 95 AND Y = 113 else
"111111111111" when X = 96 AND Y = 113 else
"111111111111" when X = 97 AND Y = 113 else
"111111111111" when X = 98 AND Y = 113 else
"111111111111" when X = 99 AND Y = 113 else
"111111111111" when X = 100 AND Y = 113 else
"111111111111" when X = 101 AND Y = 113 else
"111111111111" when X = 102 AND Y = 113 else
"111111111111" when X = 103 AND Y = 113 else
"111111111111" when X = 104 AND Y = 113 else
"111111111111" when X = 105 AND Y = 113 else
"111111111111" when X = 106 AND Y = 113 else
"111111111111" when X = 107 AND Y = 113 else
"111111111111" when X = 108 AND Y = 113 else
"111111111111" when X = 109 AND Y = 113 else
"111111111111" when X = 110 AND Y = 113 else
"111111111111" when X = 111 AND Y = 113 else
"111111111111" when X = 112 AND Y = 113 else
"111111111111" when X = 113 AND Y = 113 else
"111111111111" when X = 114 AND Y = 113 else
"111111111111" when X = 115 AND Y = 113 else
"111111111111" when X = 116 AND Y = 113 else
"111111111111" when X = 117 AND Y = 113 else
"111111111111" when X = 118 AND Y = 113 else
"111111111111" when X = 119 AND Y = 113 else
"111111111111" when X = 120 AND Y = 113 else
"111111111111" when X = 121 AND Y = 113 else
"111111111111" when X = 122 AND Y = 113 else
"111111111111" when X = 123 AND Y = 113 else
"111111111111" when X = 124 AND Y = 113 else
"111111111111" when X = 125 AND Y = 113 else
"111111111111" when X = 126 AND Y = 113 else
"111111111111" when X = 127 AND Y = 113 else
"111111111111" when X = 128 AND Y = 113 else
"111111111111" when X = 129 AND Y = 113 else
"111111111111" when X = 130 AND Y = 113 else
"111111111111" when X = 131 AND Y = 113 else
"111111111111" when X = 132 AND Y = 113 else
"111111111111" when X = 133 AND Y = 113 else
"111111111111" when X = 134 AND Y = 113 else
"111111111111" when X = 135 AND Y = 113 else
"111111111111" when X = 136 AND Y = 113 else
"111111111111" when X = 137 AND Y = 113 else
"111111111111" when X = 138 AND Y = 113 else
"111111111111" when X = 139 AND Y = 113 else
"111111111111" when X = 140 AND Y = 113 else
"111111111111" when X = 141 AND Y = 113 else
"111111111111" when X = 142 AND Y = 113 else
"111111111111" when X = 143 AND Y = 113 else
"111111111111" when X = 144 AND Y = 113 else
"111111111111" when X = 145 AND Y = 113 else
"111111111111" when X = 146 AND Y = 113 else
"111111111111" when X = 147 AND Y = 113 else
"111111111111" when X = 148 AND Y = 113 else
"111111111111" when X = 149 AND Y = 113 else
"111111111111" when X = 150 AND Y = 113 else
"111111111111" when X = 151 AND Y = 113 else
"111111111111" when X = 152 AND Y = 113 else
"111111111111" when X = 153 AND Y = 113 else
"111111111111" when X = 154 AND Y = 113 else
"111111111111" when X = 155 AND Y = 113 else
"111111111111" when X = 156 AND Y = 113 else
"111111111111" when X = 157 AND Y = 113 else
"111111111111" when X = 158 AND Y = 113 else
"111111111111" when X = 159 AND Y = 113 else
"111111111111" when X = 160 AND Y = 113 else
"111111111111" when X = 161 AND Y = 113 else
"111111111111" when X = 162 AND Y = 113 else
"111111111111" when X = 163 AND Y = 113 else
"111111111111" when X = 164 AND Y = 113 else
"111111111111" when X = 165 AND Y = 113 else
"111111111111" when X = 166 AND Y = 113 else
"111111111111" when X = 167 AND Y = 113 else
"111111111111" when X = 168 AND Y = 113 else
"111111111111" when X = 169 AND Y = 113 else
"111111111111" when X = 170 AND Y = 113 else
"111111111111" when X = 171 AND Y = 113 else
"111111111111" when X = 172 AND Y = 113 else
"111111111111" when X = 173 AND Y = 113 else
"111111111111" when X = 174 AND Y = 113 else
"111111111111" when X = 175 AND Y = 113 else
"111111111111" when X = 176 AND Y = 113 else
"111111111111" when X = 177 AND Y = 113 else
"111111111111" when X = 178 AND Y = 113 else
"111111111111" when X = 179 AND Y = 113 else
"111111111111" when X = 180 AND Y = 113 else
"111111111111" when X = 181 AND Y = 113 else
"111111111111" when X = 182 AND Y = 113 else
"111111111111" when X = 183 AND Y = 113 else
"111111111111" when X = 184 AND Y = 113 else
"111111111111" when X = 185 AND Y = 113 else
"111111111111" when X = 186 AND Y = 113 else
"111111111111" when X = 187 AND Y = 113 else
"111111111111" when X = 188 AND Y = 113 else
"111111111111" when X = 189 AND Y = 113 else
"111111111111" when X = 190 AND Y = 113 else
"111111111111" when X = 191 AND Y = 113 else
"111111111111" when X = 192 AND Y = 113 else
"111111111111" when X = 193 AND Y = 113 else
"111111111111" when X = 194 AND Y = 113 else
"111111111111" when X = 195 AND Y = 113 else
"111111111111" when X = 196 AND Y = 113 else
"111111111111" when X = 197 AND Y = 113 else
"111111111111" when X = 198 AND Y = 113 else
"111111111111" when X = 199 AND Y = 113 else
"111111111111" when X = 200 AND Y = 113 else
"111111111111" when X = 201 AND Y = 113 else
"111111111111" when X = 202 AND Y = 113 else
"111111111111" when X = 203 AND Y = 113 else
"111111111111" when X = 204 AND Y = 113 else
"111111111111" when X = 205 AND Y = 113 else
"111111111111" when X = 206 AND Y = 113 else
"111111111111" when X = 207 AND Y = 113 else
"111111111111" when X = 208 AND Y = 113 else
"111111111111" when X = 209 AND Y = 113 else
"110111011111" when X = 210 AND Y = 113 else
"110111011111" when X = 211 AND Y = 113 else
"110111011111" when X = 212 AND Y = 113 else
"110111011111" when X = 213 AND Y = 113 else
"110111011111" when X = 214 AND Y = 113 else
"110111011111" when X = 215 AND Y = 113 else
"110111011111" when X = 216 AND Y = 113 else
"110111011111" when X = 217 AND Y = 113 else
"110111011111" when X = 218 AND Y = 113 else
"110111011111" when X = 219 AND Y = 113 else
"110111011111" when X = 220 AND Y = 113 else
"110111011111" when X = 221 AND Y = 113 else
"110111011111" when X = 222 AND Y = 113 else
"110111011111" when X = 223 AND Y = 113 else
"110111011111" when X = 224 AND Y = 113 else
"110111011111" when X = 225 AND Y = 113 else
"110111011111" when X = 226 AND Y = 113 else
"110111011111" when X = 227 AND Y = 113 else
"110111011111" when X = 228 AND Y = 113 else
"110111011111" when X = 229 AND Y = 113 else
"110111011111" when X = 230 AND Y = 113 else
"110111011111" when X = 231 AND Y = 113 else
"110111011111" when X = 232 AND Y = 113 else
"110111011111" when X = 233 AND Y = 113 else
"110111011111" when X = 234 AND Y = 113 else
"110111011111" when X = 235 AND Y = 113 else
"110111011111" when X = 236 AND Y = 113 else
"110111011111" when X = 237 AND Y = 113 else
"110111011111" when X = 238 AND Y = 113 else
"110111011111" when X = 239 AND Y = 113 else
"110111011111" when X = 240 AND Y = 113 else
"110111011111" when X = 241 AND Y = 113 else
"110111011111" when X = 242 AND Y = 113 else
"110111011111" when X = 243 AND Y = 113 else
"110111011111" when X = 244 AND Y = 113 else
"110111011111" when X = 245 AND Y = 113 else
"110111011111" when X = 246 AND Y = 113 else
"110111011111" when X = 247 AND Y = 113 else
"110111011111" when X = 248 AND Y = 113 else
"110111011111" when X = 249 AND Y = 113 else
"110111011111" when X = 250 AND Y = 113 else
"110111011111" when X = 251 AND Y = 113 else
"110111011111" when X = 252 AND Y = 113 else
"110111011111" when X = 253 AND Y = 113 else
"110111011111" when X = 254 AND Y = 113 else
"110111011111" when X = 255 AND Y = 113 else
"110111011111" when X = 256 AND Y = 113 else
"110111011111" when X = 257 AND Y = 113 else
"110111011111" when X = 258 AND Y = 113 else
"110111011111" when X = 259 AND Y = 113 else
"110111011111" when X = 260 AND Y = 113 else
"110111011111" when X = 261 AND Y = 113 else
"110111011111" when X = 262 AND Y = 113 else
"110111011111" when X = 263 AND Y = 113 else
"110111011111" when X = 264 AND Y = 113 else
"110111011111" when X = 265 AND Y = 113 else
"110111011111" when X = 266 AND Y = 113 else
"110111011111" when X = 267 AND Y = 113 else
"110111011111" when X = 268 AND Y = 113 else
"110111011111" when X = 269 AND Y = 113 else
"110111011111" when X = 270 AND Y = 113 else
"110111011111" when X = 271 AND Y = 113 else
"110111011111" when X = 272 AND Y = 113 else
"110111011111" when X = 273 AND Y = 113 else
"110111011111" when X = 274 AND Y = 113 else
"110111011111" when X = 275 AND Y = 113 else
"110111011111" when X = 276 AND Y = 113 else
"110111011111" when X = 277 AND Y = 113 else
"110111011111" when X = 278 AND Y = 113 else
"110111011111" when X = 279 AND Y = 113 else
"111111111111" when X = 280 AND Y = 113 else
"111111111111" when X = 281 AND Y = 113 else
"111111111111" when X = 282 AND Y = 113 else
"111111111111" when X = 283 AND Y = 113 else
"111111111111" when X = 284 AND Y = 113 else
"111111111111" when X = 285 AND Y = 113 else
"111111111111" when X = 286 AND Y = 113 else
"111111111111" when X = 287 AND Y = 113 else
"111111111111" when X = 288 AND Y = 113 else
"111111111111" when X = 289 AND Y = 113 else
"111111111111" when X = 290 AND Y = 113 else
"111111111111" when X = 291 AND Y = 113 else
"111111111111" when X = 292 AND Y = 113 else
"111111111111" when X = 293 AND Y = 113 else
"111111111111" when X = 294 AND Y = 113 else
"111111111111" when X = 295 AND Y = 113 else
"111111111111" when X = 296 AND Y = 113 else
"111111111111" when X = 297 AND Y = 113 else
"111111111111" when X = 298 AND Y = 113 else
"111111111111" when X = 299 AND Y = 113 else
"111111111111" when X = 300 AND Y = 113 else
"111111111111" when X = 301 AND Y = 113 else
"111111111111" when X = 302 AND Y = 113 else
"111111111111" when X = 303 AND Y = 113 else
"111111111111" when X = 304 AND Y = 113 else
"110111011111" when X = 305 AND Y = 113 else
"110111011111" when X = 306 AND Y = 113 else
"110111011111" when X = 307 AND Y = 113 else
"110111011111" when X = 308 AND Y = 113 else
"110111011111" when X = 309 AND Y = 113 else
"110111011111" when X = 310 AND Y = 113 else
"110111011111" when X = 311 AND Y = 113 else
"110111011111" when X = 312 AND Y = 113 else
"110111011111" when X = 313 AND Y = 113 else
"110111011111" when X = 314 AND Y = 113 else
"110111011111" when X = 315 AND Y = 113 else
"110111011111" when X = 316 AND Y = 113 else
"110111011111" when X = 317 AND Y = 113 else
"110111011111" when X = 318 AND Y = 113 else
"110111011111" when X = 319 AND Y = 113 else
"110111011111" when X = 320 AND Y = 113 else
"110111011111" when X = 321 AND Y = 113 else
"110111011111" when X = 322 AND Y = 113 else
"110111011111" when X = 323 AND Y = 113 else
"110111011111" when X = 324 AND Y = 113 else
"100010011101" when X = 0 AND Y = 114 else
"100010011101" when X = 1 AND Y = 114 else
"100010011101" when X = 2 AND Y = 114 else
"100010011101" when X = 3 AND Y = 114 else
"100010011101" when X = 4 AND Y = 114 else
"100010011101" when X = 5 AND Y = 114 else
"100010011101" when X = 6 AND Y = 114 else
"100010011101" when X = 7 AND Y = 114 else
"100010011101" when X = 8 AND Y = 114 else
"100010011101" when X = 9 AND Y = 114 else
"100010011101" when X = 10 AND Y = 114 else
"100010011101" when X = 11 AND Y = 114 else
"100010011101" when X = 12 AND Y = 114 else
"100010011101" when X = 13 AND Y = 114 else
"100010011101" when X = 14 AND Y = 114 else
"100010011101" when X = 15 AND Y = 114 else
"100010011101" when X = 16 AND Y = 114 else
"100010011101" when X = 17 AND Y = 114 else
"100010011101" when X = 18 AND Y = 114 else
"100010011101" when X = 19 AND Y = 114 else
"100010011101" when X = 20 AND Y = 114 else
"100010011101" when X = 21 AND Y = 114 else
"100010011101" when X = 22 AND Y = 114 else
"100010011101" when X = 23 AND Y = 114 else
"100010011101" when X = 24 AND Y = 114 else
"110111011111" when X = 25 AND Y = 114 else
"110111011111" when X = 26 AND Y = 114 else
"110111011111" when X = 27 AND Y = 114 else
"110111011111" when X = 28 AND Y = 114 else
"110111011111" when X = 29 AND Y = 114 else
"110111011111" when X = 30 AND Y = 114 else
"110111011111" when X = 31 AND Y = 114 else
"110111011111" when X = 32 AND Y = 114 else
"110111011111" when X = 33 AND Y = 114 else
"110111011111" when X = 34 AND Y = 114 else
"110111011111" when X = 35 AND Y = 114 else
"110111011111" when X = 36 AND Y = 114 else
"110111011111" when X = 37 AND Y = 114 else
"110111011111" when X = 38 AND Y = 114 else
"110111011111" when X = 39 AND Y = 114 else
"110111011111" when X = 40 AND Y = 114 else
"110111011111" when X = 41 AND Y = 114 else
"110111011111" when X = 42 AND Y = 114 else
"110111011111" when X = 43 AND Y = 114 else
"110111011111" when X = 44 AND Y = 114 else
"110111011111" when X = 45 AND Y = 114 else
"110111011111" when X = 46 AND Y = 114 else
"110111011111" when X = 47 AND Y = 114 else
"110111011111" when X = 48 AND Y = 114 else
"110111011111" when X = 49 AND Y = 114 else
"110111011111" when X = 50 AND Y = 114 else
"110111011111" when X = 51 AND Y = 114 else
"110111011111" when X = 52 AND Y = 114 else
"110111011111" when X = 53 AND Y = 114 else
"110111011111" when X = 54 AND Y = 114 else
"110111011111" when X = 55 AND Y = 114 else
"110111011111" when X = 56 AND Y = 114 else
"110111011111" when X = 57 AND Y = 114 else
"110111011111" when X = 58 AND Y = 114 else
"110111011111" when X = 59 AND Y = 114 else
"110111011111" when X = 60 AND Y = 114 else
"110111011111" when X = 61 AND Y = 114 else
"110111011111" when X = 62 AND Y = 114 else
"110111011111" when X = 63 AND Y = 114 else
"110111011111" when X = 64 AND Y = 114 else
"110111011111" when X = 65 AND Y = 114 else
"110111011111" when X = 66 AND Y = 114 else
"110111011111" when X = 67 AND Y = 114 else
"110111011111" when X = 68 AND Y = 114 else
"110111011111" when X = 69 AND Y = 114 else
"111111111111" when X = 70 AND Y = 114 else
"111111111111" when X = 71 AND Y = 114 else
"111111111111" when X = 72 AND Y = 114 else
"111111111111" when X = 73 AND Y = 114 else
"111111111111" when X = 74 AND Y = 114 else
"111111111111" when X = 75 AND Y = 114 else
"111111111111" when X = 76 AND Y = 114 else
"111111111111" when X = 77 AND Y = 114 else
"111111111111" when X = 78 AND Y = 114 else
"111111111111" when X = 79 AND Y = 114 else
"111111111111" when X = 80 AND Y = 114 else
"111111111111" when X = 81 AND Y = 114 else
"111111111111" when X = 82 AND Y = 114 else
"111111111111" when X = 83 AND Y = 114 else
"111111111111" when X = 84 AND Y = 114 else
"111111111111" when X = 85 AND Y = 114 else
"111111111111" when X = 86 AND Y = 114 else
"111111111111" when X = 87 AND Y = 114 else
"111111111111" when X = 88 AND Y = 114 else
"111111111111" when X = 89 AND Y = 114 else
"111111111111" when X = 90 AND Y = 114 else
"111111111111" when X = 91 AND Y = 114 else
"111111111111" when X = 92 AND Y = 114 else
"111111111111" when X = 93 AND Y = 114 else
"111111111111" when X = 94 AND Y = 114 else
"111111111111" when X = 95 AND Y = 114 else
"111111111111" when X = 96 AND Y = 114 else
"111111111111" when X = 97 AND Y = 114 else
"111111111111" when X = 98 AND Y = 114 else
"111111111111" when X = 99 AND Y = 114 else
"111111111111" when X = 100 AND Y = 114 else
"111111111111" when X = 101 AND Y = 114 else
"111111111111" when X = 102 AND Y = 114 else
"111111111111" when X = 103 AND Y = 114 else
"111111111111" when X = 104 AND Y = 114 else
"111111111111" when X = 105 AND Y = 114 else
"111111111111" when X = 106 AND Y = 114 else
"111111111111" when X = 107 AND Y = 114 else
"111111111111" when X = 108 AND Y = 114 else
"111111111111" when X = 109 AND Y = 114 else
"111111111111" when X = 110 AND Y = 114 else
"111111111111" when X = 111 AND Y = 114 else
"111111111111" when X = 112 AND Y = 114 else
"111111111111" when X = 113 AND Y = 114 else
"111111111111" when X = 114 AND Y = 114 else
"111111111111" when X = 115 AND Y = 114 else
"111111111111" when X = 116 AND Y = 114 else
"111111111111" when X = 117 AND Y = 114 else
"111111111111" when X = 118 AND Y = 114 else
"111111111111" when X = 119 AND Y = 114 else
"111111111111" when X = 120 AND Y = 114 else
"111111111111" when X = 121 AND Y = 114 else
"111111111111" when X = 122 AND Y = 114 else
"111111111111" when X = 123 AND Y = 114 else
"111111111111" when X = 124 AND Y = 114 else
"111111111111" when X = 125 AND Y = 114 else
"111111111111" when X = 126 AND Y = 114 else
"111111111111" when X = 127 AND Y = 114 else
"111111111111" when X = 128 AND Y = 114 else
"111111111111" when X = 129 AND Y = 114 else
"111111111111" when X = 130 AND Y = 114 else
"111111111111" when X = 131 AND Y = 114 else
"111111111111" when X = 132 AND Y = 114 else
"111111111111" when X = 133 AND Y = 114 else
"111111111111" when X = 134 AND Y = 114 else
"111111111111" when X = 135 AND Y = 114 else
"111111111111" when X = 136 AND Y = 114 else
"111111111111" when X = 137 AND Y = 114 else
"111111111111" when X = 138 AND Y = 114 else
"111111111111" when X = 139 AND Y = 114 else
"111111111111" when X = 140 AND Y = 114 else
"111111111111" when X = 141 AND Y = 114 else
"111111111111" when X = 142 AND Y = 114 else
"111111111111" when X = 143 AND Y = 114 else
"111111111111" when X = 144 AND Y = 114 else
"111111111111" when X = 145 AND Y = 114 else
"111111111111" when X = 146 AND Y = 114 else
"111111111111" when X = 147 AND Y = 114 else
"111111111111" when X = 148 AND Y = 114 else
"111111111111" when X = 149 AND Y = 114 else
"111111111111" when X = 150 AND Y = 114 else
"111111111111" when X = 151 AND Y = 114 else
"111111111111" when X = 152 AND Y = 114 else
"111111111111" when X = 153 AND Y = 114 else
"111111111111" when X = 154 AND Y = 114 else
"111111111111" when X = 155 AND Y = 114 else
"111111111111" when X = 156 AND Y = 114 else
"111111111111" when X = 157 AND Y = 114 else
"111111111111" when X = 158 AND Y = 114 else
"111111111111" when X = 159 AND Y = 114 else
"111111111111" when X = 160 AND Y = 114 else
"111111111111" when X = 161 AND Y = 114 else
"111111111111" when X = 162 AND Y = 114 else
"111111111111" when X = 163 AND Y = 114 else
"111111111111" when X = 164 AND Y = 114 else
"111111111111" when X = 165 AND Y = 114 else
"111111111111" when X = 166 AND Y = 114 else
"111111111111" when X = 167 AND Y = 114 else
"111111111111" when X = 168 AND Y = 114 else
"111111111111" when X = 169 AND Y = 114 else
"111111111111" when X = 170 AND Y = 114 else
"111111111111" when X = 171 AND Y = 114 else
"111111111111" when X = 172 AND Y = 114 else
"111111111111" when X = 173 AND Y = 114 else
"111111111111" when X = 174 AND Y = 114 else
"111111111111" when X = 175 AND Y = 114 else
"111111111111" when X = 176 AND Y = 114 else
"111111111111" when X = 177 AND Y = 114 else
"111111111111" when X = 178 AND Y = 114 else
"111111111111" when X = 179 AND Y = 114 else
"111111111111" when X = 180 AND Y = 114 else
"111111111111" when X = 181 AND Y = 114 else
"111111111111" when X = 182 AND Y = 114 else
"111111111111" when X = 183 AND Y = 114 else
"111111111111" when X = 184 AND Y = 114 else
"111111111111" when X = 185 AND Y = 114 else
"111111111111" when X = 186 AND Y = 114 else
"111111111111" when X = 187 AND Y = 114 else
"111111111111" when X = 188 AND Y = 114 else
"111111111111" when X = 189 AND Y = 114 else
"111111111111" when X = 190 AND Y = 114 else
"111111111111" when X = 191 AND Y = 114 else
"111111111111" when X = 192 AND Y = 114 else
"111111111111" when X = 193 AND Y = 114 else
"111111111111" when X = 194 AND Y = 114 else
"111111111111" when X = 195 AND Y = 114 else
"111111111111" when X = 196 AND Y = 114 else
"111111111111" when X = 197 AND Y = 114 else
"111111111111" when X = 198 AND Y = 114 else
"111111111111" when X = 199 AND Y = 114 else
"111111111111" when X = 200 AND Y = 114 else
"111111111111" when X = 201 AND Y = 114 else
"111111111111" when X = 202 AND Y = 114 else
"111111111111" when X = 203 AND Y = 114 else
"111111111111" when X = 204 AND Y = 114 else
"111111111111" when X = 205 AND Y = 114 else
"111111111111" when X = 206 AND Y = 114 else
"111111111111" when X = 207 AND Y = 114 else
"111111111111" when X = 208 AND Y = 114 else
"111111111111" when X = 209 AND Y = 114 else
"110111011111" when X = 210 AND Y = 114 else
"110111011111" when X = 211 AND Y = 114 else
"110111011111" when X = 212 AND Y = 114 else
"110111011111" when X = 213 AND Y = 114 else
"110111011111" when X = 214 AND Y = 114 else
"110111011111" when X = 215 AND Y = 114 else
"110111011111" when X = 216 AND Y = 114 else
"110111011111" when X = 217 AND Y = 114 else
"110111011111" when X = 218 AND Y = 114 else
"110111011111" when X = 219 AND Y = 114 else
"110111011111" when X = 220 AND Y = 114 else
"110111011111" when X = 221 AND Y = 114 else
"110111011111" when X = 222 AND Y = 114 else
"110111011111" when X = 223 AND Y = 114 else
"110111011111" when X = 224 AND Y = 114 else
"110111011111" when X = 225 AND Y = 114 else
"110111011111" when X = 226 AND Y = 114 else
"110111011111" when X = 227 AND Y = 114 else
"110111011111" when X = 228 AND Y = 114 else
"110111011111" when X = 229 AND Y = 114 else
"110111011111" when X = 230 AND Y = 114 else
"110111011111" when X = 231 AND Y = 114 else
"110111011111" when X = 232 AND Y = 114 else
"110111011111" when X = 233 AND Y = 114 else
"110111011111" when X = 234 AND Y = 114 else
"110111011111" when X = 235 AND Y = 114 else
"110111011111" when X = 236 AND Y = 114 else
"110111011111" when X = 237 AND Y = 114 else
"110111011111" when X = 238 AND Y = 114 else
"110111011111" when X = 239 AND Y = 114 else
"110111011111" when X = 240 AND Y = 114 else
"110111011111" when X = 241 AND Y = 114 else
"110111011111" when X = 242 AND Y = 114 else
"110111011111" when X = 243 AND Y = 114 else
"110111011111" when X = 244 AND Y = 114 else
"110111011111" when X = 245 AND Y = 114 else
"110111011111" when X = 246 AND Y = 114 else
"110111011111" when X = 247 AND Y = 114 else
"110111011111" when X = 248 AND Y = 114 else
"110111011111" when X = 249 AND Y = 114 else
"110111011111" when X = 250 AND Y = 114 else
"110111011111" when X = 251 AND Y = 114 else
"110111011111" when X = 252 AND Y = 114 else
"110111011111" when X = 253 AND Y = 114 else
"110111011111" when X = 254 AND Y = 114 else
"110111011111" when X = 255 AND Y = 114 else
"110111011111" when X = 256 AND Y = 114 else
"110111011111" when X = 257 AND Y = 114 else
"110111011111" when X = 258 AND Y = 114 else
"110111011111" when X = 259 AND Y = 114 else
"110111011111" when X = 260 AND Y = 114 else
"110111011111" when X = 261 AND Y = 114 else
"110111011111" when X = 262 AND Y = 114 else
"110111011111" when X = 263 AND Y = 114 else
"110111011111" when X = 264 AND Y = 114 else
"110111011111" when X = 265 AND Y = 114 else
"110111011111" when X = 266 AND Y = 114 else
"110111011111" when X = 267 AND Y = 114 else
"110111011111" when X = 268 AND Y = 114 else
"110111011111" when X = 269 AND Y = 114 else
"110111011111" when X = 270 AND Y = 114 else
"110111011111" when X = 271 AND Y = 114 else
"110111011111" when X = 272 AND Y = 114 else
"110111011111" when X = 273 AND Y = 114 else
"110111011111" when X = 274 AND Y = 114 else
"110111011111" when X = 275 AND Y = 114 else
"110111011111" when X = 276 AND Y = 114 else
"110111011111" when X = 277 AND Y = 114 else
"110111011111" when X = 278 AND Y = 114 else
"110111011111" when X = 279 AND Y = 114 else
"111111111111" when X = 280 AND Y = 114 else
"111111111111" when X = 281 AND Y = 114 else
"111111111111" when X = 282 AND Y = 114 else
"111111111111" when X = 283 AND Y = 114 else
"111111111111" when X = 284 AND Y = 114 else
"111111111111" when X = 285 AND Y = 114 else
"111111111111" when X = 286 AND Y = 114 else
"111111111111" when X = 287 AND Y = 114 else
"111111111111" when X = 288 AND Y = 114 else
"111111111111" when X = 289 AND Y = 114 else
"111111111111" when X = 290 AND Y = 114 else
"111111111111" when X = 291 AND Y = 114 else
"111111111111" when X = 292 AND Y = 114 else
"111111111111" when X = 293 AND Y = 114 else
"111111111111" when X = 294 AND Y = 114 else
"111111111111" when X = 295 AND Y = 114 else
"111111111111" when X = 296 AND Y = 114 else
"111111111111" when X = 297 AND Y = 114 else
"111111111111" when X = 298 AND Y = 114 else
"111111111111" when X = 299 AND Y = 114 else
"111111111111" when X = 300 AND Y = 114 else
"111111111111" when X = 301 AND Y = 114 else
"111111111111" when X = 302 AND Y = 114 else
"111111111111" when X = 303 AND Y = 114 else
"111111111111" when X = 304 AND Y = 114 else
"110111011111" when X = 305 AND Y = 114 else
"110111011111" when X = 306 AND Y = 114 else
"110111011111" when X = 307 AND Y = 114 else
"110111011111" when X = 308 AND Y = 114 else
"110111011111" when X = 309 AND Y = 114 else
"110111011111" when X = 310 AND Y = 114 else
"110111011111" when X = 311 AND Y = 114 else
"110111011111" when X = 312 AND Y = 114 else
"110111011111" when X = 313 AND Y = 114 else
"110111011111" when X = 314 AND Y = 114 else
"110111011111" when X = 315 AND Y = 114 else
"110111011111" when X = 316 AND Y = 114 else
"110111011111" when X = 317 AND Y = 114 else
"110111011111" when X = 318 AND Y = 114 else
"110111011111" when X = 319 AND Y = 114 else
"110111011111" when X = 320 AND Y = 114 else
"110111011111" when X = 321 AND Y = 114 else
"110111011111" when X = 322 AND Y = 114 else
"110111011111" when X = 323 AND Y = 114 else
"110111011111" when X = 324 AND Y = 114 else
"100010011101" when X = 0 AND Y = 115 else
"100010011101" when X = 1 AND Y = 115 else
"100010011101" when X = 2 AND Y = 115 else
"100010011101" when X = 3 AND Y = 115 else
"100010011101" when X = 4 AND Y = 115 else
"100010011101" when X = 5 AND Y = 115 else
"100010011101" when X = 6 AND Y = 115 else
"100010011101" when X = 7 AND Y = 115 else
"100010011101" when X = 8 AND Y = 115 else
"100010011101" when X = 9 AND Y = 115 else
"100010011101" when X = 10 AND Y = 115 else
"100010011101" when X = 11 AND Y = 115 else
"100010011101" when X = 12 AND Y = 115 else
"100010011101" when X = 13 AND Y = 115 else
"100010011101" when X = 14 AND Y = 115 else
"100010011101" when X = 15 AND Y = 115 else
"100010011101" when X = 16 AND Y = 115 else
"100010011101" when X = 17 AND Y = 115 else
"100010011101" when X = 18 AND Y = 115 else
"100010011101" when X = 19 AND Y = 115 else
"100010011101" when X = 20 AND Y = 115 else
"100010011101" when X = 21 AND Y = 115 else
"100010011101" when X = 22 AND Y = 115 else
"100010011101" when X = 23 AND Y = 115 else
"100010011101" when X = 24 AND Y = 115 else
"100010011101" when X = 25 AND Y = 115 else
"100010011101" when X = 26 AND Y = 115 else
"100010011101" when X = 27 AND Y = 115 else
"100010011101" when X = 28 AND Y = 115 else
"100010011101" when X = 29 AND Y = 115 else
"110111011111" when X = 30 AND Y = 115 else
"110111011111" when X = 31 AND Y = 115 else
"110111011111" when X = 32 AND Y = 115 else
"110111011111" when X = 33 AND Y = 115 else
"110111011111" when X = 34 AND Y = 115 else
"110111011111" when X = 35 AND Y = 115 else
"110111011111" when X = 36 AND Y = 115 else
"110111011111" when X = 37 AND Y = 115 else
"110111011111" when X = 38 AND Y = 115 else
"110111011111" when X = 39 AND Y = 115 else
"110111011111" when X = 40 AND Y = 115 else
"110111011111" when X = 41 AND Y = 115 else
"110111011111" when X = 42 AND Y = 115 else
"110111011111" when X = 43 AND Y = 115 else
"110111011111" when X = 44 AND Y = 115 else
"110111011111" when X = 45 AND Y = 115 else
"110111011111" when X = 46 AND Y = 115 else
"110111011111" when X = 47 AND Y = 115 else
"110111011111" when X = 48 AND Y = 115 else
"110111011111" when X = 49 AND Y = 115 else
"110111011111" when X = 50 AND Y = 115 else
"110111011111" when X = 51 AND Y = 115 else
"110111011111" when X = 52 AND Y = 115 else
"110111011111" when X = 53 AND Y = 115 else
"110111011111" when X = 54 AND Y = 115 else
"110111011111" when X = 55 AND Y = 115 else
"110111011111" when X = 56 AND Y = 115 else
"110111011111" when X = 57 AND Y = 115 else
"110111011111" when X = 58 AND Y = 115 else
"110111011111" when X = 59 AND Y = 115 else
"110111011111" when X = 60 AND Y = 115 else
"110111011111" when X = 61 AND Y = 115 else
"110111011111" when X = 62 AND Y = 115 else
"110111011111" when X = 63 AND Y = 115 else
"110111011111" when X = 64 AND Y = 115 else
"110111011111" when X = 65 AND Y = 115 else
"110111011111" when X = 66 AND Y = 115 else
"110111011111" when X = 67 AND Y = 115 else
"110111011111" when X = 68 AND Y = 115 else
"110111011111" when X = 69 AND Y = 115 else
"110111011111" when X = 70 AND Y = 115 else
"110111011111" when X = 71 AND Y = 115 else
"110111011111" when X = 72 AND Y = 115 else
"110111011111" when X = 73 AND Y = 115 else
"110111011111" when X = 74 AND Y = 115 else
"110111011111" when X = 75 AND Y = 115 else
"110111011111" when X = 76 AND Y = 115 else
"110111011111" when X = 77 AND Y = 115 else
"110111011111" when X = 78 AND Y = 115 else
"110111011111" when X = 79 AND Y = 115 else
"110111011111" when X = 80 AND Y = 115 else
"110111011111" when X = 81 AND Y = 115 else
"110111011111" when X = 82 AND Y = 115 else
"110111011111" when X = 83 AND Y = 115 else
"110111011111" when X = 84 AND Y = 115 else
"110111011111" when X = 85 AND Y = 115 else
"110111011111" when X = 86 AND Y = 115 else
"110111011111" when X = 87 AND Y = 115 else
"110111011111" when X = 88 AND Y = 115 else
"110111011111" when X = 89 AND Y = 115 else
"110111011111" when X = 90 AND Y = 115 else
"110111011111" when X = 91 AND Y = 115 else
"110111011111" when X = 92 AND Y = 115 else
"110111011111" when X = 93 AND Y = 115 else
"110111011111" when X = 94 AND Y = 115 else
"110111011111" when X = 95 AND Y = 115 else
"110111011111" when X = 96 AND Y = 115 else
"110111011111" when X = 97 AND Y = 115 else
"110111011111" when X = 98 AND Y = 115 else
"110111011111" when X = 99 AND Y = 115 else
"110111011111" when X = 100 AND Y = 115 else
"110111011111" when X = 101 AND Y = 115 else
"110111011111" when X = 102 AND Y = 115 else
"110111011111" when X = 103 AND Y = 115 else
"110111011111" when X = 104 AND Y = 115 else
"110111011111" when X = 105 AND Y = 115 else
"110111011111" when X = 106 AND Y = 115 else
"110111011111" when X = 107 AND Y = 115 else
"110111011111" when X = 108 AND Y = 115 else
"110111011111" when X = 109 AND Y = 115 else
"110111011111" when X = 110 AND Y = 115 else
"110111011111" when X = 111 AND Y = 115 else
"110111011111" when X = 112 AND Y = 115 else
"110111011111" when X = 113 AND Y = 115 else
"110111011111" when X = 114 AND Y = 115 else
"110111011111" when X = 115 AND Y = 115 else
"110111011111" when X = 116 AND Y = 115 else
"110111011111" when X = 117 AND Y = 115 else
"110111011111" when X = 118 AND Y = 115 else
"110111011111" when X = 119 AND Y = 115 else
"110111011111" when X = 120 AND Y = 115 else
"110111011111" when X = 121 AND Y = 115 else
"110111011111" when X = 122 AND Y = 115 else
"110111011111" when X = 123 AND Y = 115 else
"110111011111" when X = 124 AND Y = 115 else
"110111011111" when X = 125 AND Y = 115 else
"110111011111" when X = 126 AND Y = 115 else
"110111011111" when X = 127 AND Y = 115 else
"110111011111" when X = 128 AND Y = 115 else
"110111011111" when X = 129 AND Y = 115 else
"110111011111" when X = 130 AND Y = 115 else
"110111011111" when X = 131 AND Y = 115 else
"110111011111" when X = 132 AND Y = 115 else
"110111011111" when X = 133 AND Y = 115 else
"110111011111" when X = 134 AND Y = 115 else
"110111011111" when X = 135 AND Y = 115 else
"110111011111" when X = 136 AND Y = 115 else
"110111011111" when X = 137 AND Y = 115 else
"110111011111" when X = 138 AND Y = 115 else
"110111011111" when X = 139 AND Y = 115 else
"110111011111" when X = 140 AND Y = 115 else
"110111011111" when X = 141 AND Y = 115 else
"110111011111" when X = 142 AND Y = 115 else
"110111011111" when X = 143 AND Y = 115 else
"110111011111" when X = 144 AND Y = 115 else
"111111111111" when X = 145 AND Y = 115 else
"111111111111" when X = 146 AND Y = 115 else
"111111111111" when X = 147 AND Y = 115 else
"111111111111" when X = 148 AND Y = 115 else
"111111111111" when X = 149 AND Y = 115 else
"111111111111" when X = 150 AND Y = 115 else
"111111111111" when X = 151 AND Y = 115 else
"111111111111" when X = 152 AND Y = 115 else
"111111111111" when X = 153 AND Y = 115 else
"111111111111" when X = 154 AND Y = 115 else
"111111111111" when X = 155 AND Y = 115 else
"111111111111" when X = 156 AND Y = 115 else
"111111111111" when X = 157 AND Y = 115 else
"111111111111" when X = 158 AND Y = 115 else
"111111111111" when X = 159 AND Y = 115 else
"111111111111" when X = 160 AND Y = 115 else
"111111111111" when X = 161 AND Y = 115 else
"111111111111" when X = 162 AND Y = 115 else
"111111111111" when X = 163 AND Y = 115 else
"111111111111" when X = 164 AND Y = 115 else
"111111111111" when X = 165 AND Y = 115 else
"111111111111" when X = 166 AND Y = 115 else
"111111111111" when X = 167 AND Y = 115 else
"111111111111" when X = 168 AND Y = 115 else
"111111111111" when X = 169 AND Y = 115 else
"111111111111" when X = 170 AND Y = 115 else
"111111111111" when X = 171 AND Y = 115 else
"111111111111" when X = 172 AND Y = 115 else
"111111111111" when X = 173 AND Y = 115 else
"111111111111" when X = 174 AND Y = 115 else
"111111111111" when X = 175 AND Y = 115 else
"111111111111" when X = 176 AND Y = 115 else
"111111111111" when X = 177 AND Y = 115 else
"111111111111" when X = 178 AND Y = 115 else
"111111111111" when X = 179 AND Y = 115 else
"111111111111" when X = 180 AND Y = 115 else
"111111111111" when X = 181 AND Y = 115 else
"111111111111" when X = 182 AND Y = 115 else
"111111111111" when X = 183 AND Y = 115 else
"111111111111" when X = 184 AND Y = 115 else
"111111111111" when X = 185 AND Y = 115 else
"111111111111" when X = 186 AND Y = 115 else
"111111111111" when X = 187 AND Y = 115 else
"111111111111" when X = 188 AND Y = 115 else
"111111111111" when X = 189 AND Y = 115 else
"111111111111" when X = 190 AND Y = 115 else
"111111111111" when X = 191 AND Y = 115 else
"111111111111" when X = 192 AND Y = 115 else
"111111111111" when X = 193 AND Y = 115 else
"111111111111" when X = 194 AND Y = 115 else
"111111111111" when X = 195 AND Y = 115 else
"111111111111" when X = 196 AND Y = 115 else
"111111111111" when X = 197 AND Y = 115 else
"111111111111" when X = 198 AND Y = 115 else
"111111111111" when X = 199 AND Y = 115 else
"111111111111" when X = 200 AND Y = 115 else
"111111111111" when X = 201 AND Y = 115 else
"111111111111" when X = 202 AND Y = 115 else
"111111111111" when X = 203 AND Y = 115 else
"111111111111" when X = 204 AND Y = 115 else
"110111011111" when X = 205 AND Y = 115 else
"110111011111" when X = 206 AND Y = 115 else
"110111011111" when X = 207 AND Y = 115 else
"110111011111" when X = 208 AND Y = 115 else
"110111011111" when X = 209 AND Y = 115 else
"110111011111" when X = 210 AND Y = 115 else
"110111011111" when X = 211 AND Y = 115 else
"110111011111" when X = 212 AND Y = 115 else
"110111011111" when X = 213 AND Y = 115 else
"110111011111" when X = 214 AND Y = 115 else
"110111011111" when X = 215 AND Y = 115 else
"110111011111" when X = 216 AND Y = 115 else
"110111011111" when X = 217 AND Y = 115 else
"110111011111" when X = 218 AND Y = 115 else
"110111011111" when X = 219 AND Y = 115 else
"110111011111" when X = 220 AND Y = 115 else
"110111011111" when X = 221 AND Y = 115 else
"110111011111" when X = 222 AND Y = 115 else
"110111011111" when X = 223 AND Y = 115 else
"110111011111" when X = 224 AND Y = 115 else
"110111011111" when X = 225 AND Y = 115 else
"110111011111" when X = 226 AND Y = 115 else
"110111011111" when X = 227 AND Y = 115 else
"110111011111" when X = 228 AND Y = 115 else
"110111011111" when X = 229 AND Y = 115 else
"110111011111" when X = 230 AND Y = 115 else
"110111011111" when X = 231 AND Y = 115 else
"110111011111" when X = 232 AND Y = 115 else
"110111011111" when X = 233 AND Y = 115 else
"110111011111" when X = 234 AND Y = 115 else
"110111011111" when X = 235 AND Y = 115 else
"110111011111" when X = 236 AND Y = 115 else
"110111011111" when X = 237 AND Y = 115 else
"110111011111" when X = 238 AND Y = 115 else
"110111011111" when X = 239 AND Y = 115 else
"110111011111" when X = 240 AND Y = 115 else
"110111011111" when X = 241 AND Y = 115 else
"110111011111" when X = 242 AND Y = 115 else
"110111011111" when X = 243 AND Y = 115 else
"110111011111" when X = 244 AND Y = 115 else
"110111011111" when X = 245 AND Y = 115 else
"110111011111" when X = 246 AND Y = 115 else
"110111011111" when X = 247 AND Y = 115 else
"110111011111" when X = 248 AND Y = 115 else
"110111011111" when X = 249 AND Y = 115 else
"110111011111" when X = 250 AND Y = 115 else
"110111011111" when X = 251 AND Y = 115 else
"110111011111" when X = 252 AND Y = 115 else
"110111011111" when X = 253 AND Y = 115 else
"110111011111" when X = 254 AND Y = 115 else
"110111011111" when X = 255 AND Y = 115 else
"110111011111" when X = 256 AND Y = 115 else
"110111011111" when X = 257 AND Y = 115 else
"110111011111" when X = 258 AND Y = 115 else
"110111011111" when X = 259 AND Y = 115 else
"110111011111" when X = 260 AND Y = 115 else
"110111011111" when X = 261 AND Y = 115 else
"110111011111" when X = 262 AND Y = 115 else
"110111011111" when X = 263 AND Y = 115 else
"110111011111" when X = 264 AND Y = 115 else
"110111011111" when X = 265 AND Y = 115 else
"110111011111" when X = 266 AND Y = 115 else
"110111011111" when X = 267 AND Y = 115 else
"110111011111" when X = 268 AND Y = 115 else
"110111011111" when X = 269 AND Y = 115 else
"110111011111" when X = 270 AND Y = 115 else
"110111011111" when X = 271 AND Y = 115 else
"110111011111" when X = 272 AND Y = 115 else
"110111011111" when X = 273 AND Y = 115 else
"110111011111" when X = 274 AND Y = 115 else
"110111011111" when X = 275 AND Y = 115 else
"110111011111" when X = 276 AND Y = 115 else
"110111011111" when X = 277 AND Y = 115 else
"110111011111" when X = 278 AND Y = 115 else
"110111011111" when X = 279 AND Y = 115 else
"111111111111" when X = 280 AND Y = 115 else
"111111111111" when X = 281 AND Y = 115 else
"111111111111" when X = 282 AND Y = 115 else
"111111111111" when X = 283 AND Y = 115 else
"111111111111" when X = 284 AND Y = 115 else
"111111111111" when X = 285 AND Y = 115 else
"111111111111" when X = 286 AND Y = 115 else
"111111111111" when X = 287 AND Y = 115 else
"111111111111" when X = 288 AND Y = 115 else
"111111111111" when X = 289 AND Y = 115 else
"111111111111" when X = 290 AND Y = 115 else
"111111111111" when X = 291 AND Y = 115 else
"111111111111" when X = 292 AND Y = 115 else
"111111111111" when X = 293 AND Y = 115 else
"111111111111" when X = 294 AND Y = 115 else
"111111111111" when X = 295 AND Y = 115 else
"111111111111" when X = 296 AND Y = 115 else
"111111111111" when X = 297 AND Y = 115 else
"111111111111" when X = 298 AND Y = 115 else
"111111111111" when X = 299 AND Y = 115 else
"110111011111" when X = 300 AND Y = 115 else
"110111011111" when X = 301 AND Y = 115 else
"110111011111" when X = 302 AND Y = 115 else
"110111011111" when X = 303 AND Y = 115 else
"110111011111" when X = 304 AND Y = 115 else
"110111011111" when X = 305 AND Y = 115 else
"110111011111" when X = 306 AND Y = 115 else
"110111011111" when X = 307 AND Y = 115 else
"110111011111" when X = 308 AND Y = 115 else
"110111011111" when X = 309 AND Y = 115 else
"110111011111" when X = 310 AND Y = 115 else
"110111011111" when X = 311 AND Y = 115 else
"110111011111" when X = 312 AND Y = 115 else
"110111011111" when X = 313 AND Y = 115 else
"110111011111" when X = 314 AND Y = 115 else
"110111011111" when X = 315 AND Y = 115 else
"110111011111" when X = 316 AND Y = 115 else
"110111011111" when X = 317 AND Y = 115 else
"110111011111" when X = 318 AND Y = 115 else
"110111011111" when X = 319 AND Y = 115 else
"110111011111" when X = 320 AND Y = 115 else
"110111011111" when X = 321 AND Y = 115 else
"110111011111" when X = 322 AND Y = 115 else
"110111011111" when X = 323 AND Y = 115 else
"110111011111" when X = 324 AND Y = 115 else
"100010011101" when X = 0 AND Y = 116 else
"100010011101" when X = 1 AND Y = 116 else
"100010011101" when X = 2 AND Y = 116 else
"100010011101" when X = 3 AND Y = 116 else
"100010011101" when X = 4 AND Y = 116 else
"100010011101" when X = 5 AND Y = 116 else
"100010011101" when X = 6 AND Y = 116 else
"100010011101" when X = 7 AND Y = 116 else
"100010011101" when X = 8 AND Y = 116 else
"100010011101" when X = 9 AND Y = 116 else
"100010011101" when X = 10 AND Y = 116 else
"100010011101" when X = 11 AND Y = 116 else
"100010011101" when X = 12 AND Y = 116 else
"100010011101" when X = 13 AND Y = 116 else
"100010011101" when X = 14 AND Y = 116 else
"100010011101" when X = 15 AND Y = 116 else
"100010011101" when X = 16 AND Y = 116 else
"100010011101" when X = 17 AND Y = 116 else
"100010011101" when X = 18 AND Y = 116 else
"100010011101" when X = 19 AND Y = 116 else
"100010011101" when X = 20 AND Y = 116 else
"100010011101" when X = 21 AND Y = 116 else
"100010011101" when X = 22 AND Y = 116 else
"100010011101" when X = 23 AND Y = 116 else
"100010011101" when X = 24 AND Y = 116 else
"100010011101" when X = 25 AND Y = 116 else
"100010011101" when X = 26 AND Y = 116 else
"100010011101" when X = 27 AND Y = 116 else
"100010011101" when X = 28 AND Y = 116 else
"100010011101" when X = 29 AND Y = 116 else
"110111011111" when X = 30 AND Y = 116 else
"110111011111" when X = 31 AND Y = 116 else
"110111011111" when X = 32 AND Y = 116 else
"110111011111" when X = 33 AND Y = 116 else
"110111011111" when X = 34 AND Y = 116 else
"110111011111" when X = 35 AND Y = 116 else
"110111011111" when X = 36 AND Y = 116 else
"110111011111" when X = 37 AND Y = 116 else
"110111011111" when X = 38 AND Y = 116 else
"110111011111" when X = 39 AND Y = 116 else
"110111011111" when X = 40 AND Y = 116 else
"110111011111" when X = 41 AND Y = 116 else
"110111011111" when X = 42 AND Y = 116 else
"110111011111" when X = 43 AND Y = 116 else
"110111011111" when X = 44 AND Y = 116 else
"110111011111" when X = 45 AND Y = 116 else
"110111011111" when X = 46 AND Y = 116 else
"110111011111" when X = 47 AND Y = 116 else
"110111011111" when X = 48 AND Y = 116 else
"110111011111" when X = 49 AND Y = 116 else
"110111011111" when X = 50 AND Y = 116 else
"110111011111" when X = 51 AND Y = 116 else
"110111011111" when X = 52 AND Y = 116 else
"110111011111" when X = 53 AND Y = 116 else
"110111011111" when X = 54 AND Y = 116 else
"110111011111" when X = 55 AND Y = 116 else
"110111011111" when X = 56 AND Y = 116 else
"110111011111" when X = 57 AND Y = 116 else
"110111011111" when X = 58 AND Y = 116 else
"110111011111" when X = 59 AND Y = 116 else
"110111011111" when X = 60 AND Y = 116 else
"110111011111" when X = 61 AND Y = 116 else
"110111011111" when X = 62 AND Y = 116 else
"110111011111" when X = 63 AND Y = 116 else
"110111011111" when X = 64 AND Y = 116 else
"110111011111" when X = 65 AND Y = 116 else
"110111011111" when X = 66 AND Y = 116 else
"110111011111" when X = 67 AND Y = 116 else
"110111011111" when X = 68 AND Y = 116 else
"110111011111" when X = 69 AND Y = 116 else
"110111011111" when X = 70 AND Y = 116 else
"110111011111" when X = 71 AND Y = 116 else
"110111011111" when X = 72 AND Y = 116 else
"110111011111" when X = 73 AND Y = 116 else
"110111011111" when X = 74 AND Y = 116 else
"110111011111" when X = 75 AND Y = 116 else
"110111011111" when X = 76 AND Y = 116 else
"110111011111" when X = 77 AND Y = 116 else
"110111011111" when X = 78 AND Y = 116 else
"110111011111" when X = 79 AND Y = 116 else
"110111011111" when X = 80 AND Y = 116 else
"110111011111" when X = 81 AND Y = 116 else
"110111011111" when X = 82 AND Y = 116 else
"110111011111" when X = 83 AND Y = 116 else
"110111011111" when X = 84 AND Y = 116 else
"110111011111" when X = 85 AND Y = 116 else
"110111011111" when X = 86 AND Y = 116 else
"110111011111" when X = 87 AND Y = 116 else
"110111011111" when X = 88 AND Y = 116 else
"110111011111" when X = 89 AND Y = 116 else
"110111011111" when X = 90 AND Y = 116 else
"110111011111" when X = 91 AND Y = 116 else
"110111011111" when X = 92 AND Y = 116 else
"110111011111" when X = 93 AND Y = 116 else
"110111011111" when X = 94 AND Y = 116 else
"110111011111" when X = 95 AND Y = 116 else
"110111011111" when X = 96 AND Y = 116 else
"110111011111" when X = 97 AND Y = 116 else
"110111011111" when X = 98 AND Y = 116 else
"110111011111" when X = 99 AND Y = 116 else
"110111011111" when X = 100 AND Y = 116 else
"110111011111" when X = 101 AND Y = 116 else
"110111011111" when X = 102 AND Y = 116 else
"110111011111" when X = 103 AND Y = 116 else
"110111011111" when X = 104 AND Y = 116 else
"110111011111" when X = 105 AND Y = 116 else
"110111011111" when X = 106 AND Y = 116 else
"110111011111" when X = 107 AND Y = 116 else
"110111011111" when X = 108 AND Y = 116 else
"110111011111" when X = 109 AND Y = 116 else
"110111011111" when X = 110 AND Y = 116 else
"110111011111" when X = 111 AND Y = 116 else
"110111011111" when X = 112 AND Y = 116 else
"110111011111" when X = 113 AND Y = 116 else
"110111011111" when X = 114 AND Y = 116 else
"110111011111" when X = 115 AND Y = 116 else
"110111011111" when X = 116 AND Y = 116 else
"110111011111" when X = 117 AND Y = 116 else
"110111011111" when X = 118 AND Y = 116 else
"110111011111" when X = 119 AND Y = 116 else
"110111011111" when X = 120 AND Y = 116 else
"110111011111" when X = 121 AND Y = 116 else
"110111011111" when X = 122 AND Y = 116 else
"110111011111" when X = 123 AND Y = 116 else
"110111011111" when X = 124 AND Y = 116 else
"110111011111" when X = 125 AND Y = 116 else
"110111011111" when X = 126 AND Y = 116 else
"110111011111" when X = 127 AND Y = 116 else
"110111011111" when X = 128 AND Y = 116 else
"110111011111" when X = 129 AND Y = 116 else
"110111011111" when X = 130 AND Y = 116 else
"110111011111" when X = 131 AND Y = 116 else
"110111011111" when X = 132 AND Y = 116 else
"110111011111" when X = 133 AND Y = 116 else
"110111011111" when X = 134 AND Y = 116 else
"110111011111" when X = 135 AND Y = 116 else
"110111011111" when X = 136 AND Y = 116 else
"110111011111" when X = 137 AND Y = 116 else
"110111011111" when X = 138 AND Y = 116 else
"110111011111" when X = 139 AND Y = 116 else
"110111011111" when X = 140 AND Y = 116 else
"110111011111" when X = 141 AND Y = 116 else
"110111011111" when X = 142 AND Y = 116 else
"110111011111" when X = 143 AND Y = 116 else
"110111011111" when X = 144 AND Y = 116 else
"111111111111" when X = 145 AND Y = 116 else
"111111111111" when X = 146 AND Y = 116 else
"111111111111" when X = 147 AND Y = 116 else
"111111111111" when X = 148 AND Y = 116 else
"111111111111" when X = 149 AND Y = 116 else
"111111111111" when X = 150 AND Y = 116 else
"111111111111" when X = 151 AND Y = 116 else
"111111111111" when X = 152 AND Y = 116 else
"111111111111" when X = 153 AND Y = 116 else
"111111111111" when X = 154 AND Y = 116 else
"111111111111" when X = 155 AND Y = 116 else
"111111111111" when X = 156 AND Y = 116 else
"111111111111" when X = 157 AND Y = 116 else
"111111111111" when X = 158 AND Y = 116 else
"111111111111" when X = 159 AND Y = 116 else
"111111111111" when X = 160 AND Y = 116 else
"111111111111" when X = 161 AND Y = 116 else
"111111111111" when X = 162 AND Y = 116 else
"111111111111" when X = 163 AND Y = 116 else
"111111111111" when X = 164 AND Y = 116 else
"111111111111" when X = 165 AND Y = 116 else
"111111111111" when X = 166 AND Y = 116 else
"111111111111" when X = 167 AND Y = 116 else
"111111111111" when X = 168 AND Y = 116 else
"111111111111" when X = 169 AND Y = 116 else
"111111111111" when X = 170 AND Y = 116 else
"111111111111" when X = 171 AND Y = 116 else
"111111111111" when X = 172 AND Y = 116 else
"111111111111" when X = 173 AND Y = 116 else
"111111111111" when X = 174 AND Y = 116 else
"111111111111" when X = 175 AND Y = 116 else
"111111111111" when X = 176 AND Y = 116 else
"111111111111" when X = 177 AND Y = 116 else
"111111111111" when X = 178 AND Y = 116 else
"111111111111" when X = 179 AND Y = 116 else
"111111111111" when X = 180 AND Y = 116 else
"111111111111" when X = 181 AND Y = 116 else
"111111111111" when X = 182 AND Y = 116 else
"111111111111" when X = 183 AND Y = 116 else
"111111111111" when X = 184 AND Y = 116 else
"111111111111" when X = 185 AND Y = 116 else
"111111111111" when X = 186 AND Y = 116 else
"111111111111" when X = 187 AND Y = 116 else
"111111111111" when X = 188 AND Y = 116 else
"111111111111" when X = 189 AND Y = 116 else
"111111111111" when X = 190 AND Y = 116 else
"111111111111" when X = 191 AND Y = 116 else
"111111111111" when X = 192 AND Y = 116 else
"111111111111" when X = 193 AND Y = 116 else
"111111111111" when X = 194 AND Y = 116 else
"111111111111" when X = 195 AND Y = 116 else
"111111111111" when X = 196 AND Y = 116 else
"111111111111" when X = 197 AND Y = 116 else
"111111111111" when X = 198 AND Y = 116 else
"111111111111" when X = 199 AND Y = 116 else
"111111111111" when X = 200 AND Y = 116 else
"111111111111" when X = 201 AND Y = 116 else
"111111111111" when X = 202 AND Y = 116 else
"111111111111" when X = 203 AND Y = 116 else
"111111111111" when X = 204 AND Y = 116 else
"110111011111" when X = 205 AND Y = 116 else
"110111011111" when X = 206 AND Y = 116 else
"110111011111" when X = 207 AND Y = 116 else
"110111011111" when X = 208 AND Y = 116 else
"110111011111" when X = 209 AND Y = 116 else
"110111011111" when X = 210 AND Y = 116 else
"110111011111" when X = 211 AND Y = 116 else
"110111011111" when X = 212 AND Y = 116 else
"110111011111" when X = 213 AND Y = 116 else
"110111011111" when X = 214 AND Y = 116 else
"110111011111" when X = 215 AND Y = 116 else
"110111011111" when X = 216 AND Y = 116 else
"110111011111" when X = 217 AND Y = 116 else
"110111011111" when X = 218 AND Y = 116 else
"110111011111" when X = 219 AND Y = 116 else
"110111011111" when X = 220 AND Y = 116 else
"110111011111" when X = 221 AND Y = 116 else
"110111011111" when X = 222 AND Y = 116 else
"110111011111" when X = 223 AND Y = 116 else
"110111011111" when X = 224 AND Y = 116 else
"110111011111" when X = 225 AND Y = 116 else
"110111011111" when X = 226 AND Y = 116 else
"110111011111" when X = 227 AND Y = 116 else
"110111011111" when X = 228 AND Y = 116 else
"110111011111" when X = 229 AND Y = 116 else
"110111011111" when X = 230 AND Y = 116 else
"110111011111" when X = 231 AND Y = 116 else
"110111011111" when X = 232 AND Y = 116 else
"110111011111" when X = 233 AND Y = 116 else
"110111011111" when X = 234 AND Y = 116 else
"110111011111" when X = 235 AND Y = 116 else
"110111011111" when X = 236 AND Y = 116 else
"110111011111" when X = 237 AND Y = 116 else
"110111011111" when X = 238 AND Y = 116 else
"110111011111" when X = 239 AND Y = 116 else
"110111011111" when X = 240 AND Y = 116 else
"110111011111" when X = 241 AND Y = 116 else
"110111011111" when X = 242 AND Y = 116 else
"110111011111" when X = 243 AND Y = 116 else
"110111011111" when X = 244 AND Y = 116 else
"110111011111" when X = 245 AND Y = 116 else
"110111011111" when X = 246 AND Y = 116 else
"110111011111" when X = 247 AND Y = 116 else
"110111011111" when X = 248 AND Y = 116 else
"110111011111" when X = 249 AND Y = 116 else
"110111011111" when X = 250 AND Y = 116 else
"110111011111" when X = 251 AND Y = 116 else
"110111011111" when X = 252 AND Y = 116 else
"110111011111" when X = 253 AND Y = 116 else
"110111011111" when X = 254 AND Y = 116 else
"110111011111" when X = 255 AND Y = 116 else
"110111011111" when X = 256 AND Y = 116 else
"110111011111" when X = 257 AND Y = 116 else
"110111011111" when X = 258 AND Y = 116 else
"110111011111" when X = 259 AND Y = 116 else
"110111011111" when X = 260 AND Y = 116 else
"110111011111" when X = 261 AND Y = 116 else
"110111011111" when X = 262 AND Y = 116 else
"110111011111" when X = 263 AND Y = 116 else
"110111011111" when X = 264 AND Y = 116 else
"110111011111" when X = 265 AND Y = 116 else
"110111011111" when X = 266 AND Y = 116 else
"110111011111" when X = 267 AND Y = 116 else
"110111011111" when X = 268 AND Y = 116 else
"110111011111" when X = 269 AND Y = 116 else
"110111011111" when X = 270 AND Y = 116 else
"110111011111" when X = 271 AND Y = 116 else
"110111011111" when X = 272 AND Y = 116 else
"110111011111" when X = 273 AND Y = 116 else
"110111011111" when X = 274 AND Y = 116 else
"110111011111" when X = 275 AND Y = 116 else
"110111011111" when X = 276 AND Y = 116 else
"110111011111" when X = 277 AND Y = 116 else
"110111011111" when X = 278 AND Y = 116 else
"110111011111" when X = 279 AND Y = 116 else
"111111111111" when X = 280 AND Y = 116 else
"111111111111" when X = 281 AND Y = 116 else
"111111111111" when X = 282 AND Y = 116 else
"111111111111" when X = 283 AND Y = 116 else
"111111111111" when X = 284 AND Y = 116 else
"111111111111" when X = 285 AND Y = 116 else
"111111111111" when X = 286 AND Y = 116 else
"111111111111" when X = 287 AND Y = 116 else
"111111111111" when X = 288 AND Y = 116 else
"111111111111" when X = 289 AND Y = 116 else
"111111111111" when X = 290 AND Y = 116 else
"111111111111" when X = 291 AND Y = 116 else
"111111111111" when X = 292 AND Y = 116 else
"111111111111" when X = 293 AND Y = 116 else
"111111111111" when X = 294 AND Y = 116 else
"111111111111" when X = 295 AND Y = 116 else
"111111111111" when X = 296 AND Y = 116 else
"111111111111" when X = 297 AND Y = 116 else
"111111111111" when X = 298 AND Y = 116 else
"111111111111" when X = 299 AND Y = 116 else
"110111011111" when X = 300 AND Y = 116 else
"110111011111" when X = 301 AND Y = 116 else
"110111011111" when X = 302 AND Y = 116 else
"110111011111" when X = 303 AND Y = 116 else
"110111011111" when X = 304 AND Y = 116 else
"110111011111" when X = 305 AND Y = 116 else
"110111011111" when X = 306 AND Y = 116 else
"110111011111" when X = 307 AND Y = 116 else
"110111011111" when X = 308 AND Y = 116 else
"110111011111" when X = 309 AND Y = 116 else
"110111011111" when X = 310 AND Y = 116 else
"110111011111" when X = 311 AND Y = 116 else
"110111011111" when X = 312 AND Y = 116 else
"110111011111" when X = 313 AND Y = 116 else
"110111011111" when X = 314 AND Y = 116 else
"110111011111" when X = 315 AND Y = 116 else
"110111011111" when X = 316 AND Y = 116 else
"110111011111" when X = 317 AND Y = 116 else
"110111011111" when X = 318 AND Y = 116 else
"110111011111" when X = 319 AND Y = 116 else
"110111011111" when X = 320 AND Y = 116 else
"110111011111" when X = 321 AND Y = 116 else
"110111011111" when X = 322 AND Y = 116 else
"110111011111" when X = 323 AND Y = 116 else
"110111011111" when X = 324 AND Y = 116 else
"100010011101" when X = 0 AND Y = 117 else
"100010011101" when X = 1 AND Y = 117 else
"100010011101" when X = 2 AND Y = 117 else
"100010011101" when X = 3 AND Y = 117 else
"100010011101" when X = 4 AND Y = 117 else
"100010011101" when X = 5 AND Y = 117 else
"100010011101" when X = 6 AND Y = 117 else
"100010011101" when X = 7 AND Y = 117 else
"100010011101" when X = 8 AND Y = 117 else
"100010011101" when X = 9 AND Y = 117 else
"100010011101" when X = 10 AND Y = 117 else
"100010011101" when X = 11 AND Y = 117 else
"100010011101" when X = 12 AND Y = 117 else
"100010011101" when X = 13 AND Y = 117 else
"100010011101" when X = 14 AND Y = 117 else
"100010011101" when X = 15 AND Y = 117 else
"100010011101" when X = 16 AND Y = 117 else
"100010011101" when X = 17 AND Y = 117 else
"100010011101" when X = 18 AND Y = 117 else
"100010011101" when X = 19 AND Y = 117 else
"100010011101" when X = 20 AND Y = 117 else
"100010011101" when X = 21 AND Y = 117 else
"100010011101" when X = 22 AND Y = 117 else
"100010011101" when X = 23 AND Y = 117 else
"100010011101" when X = 24 AND Y = 117 else
"100010011101" when X = 25 AND Y = 117 else
"100010011101" when X = 26 AND Y = 117 else
"100010011101" when X = 27 AND Y = 117 else
"100010011101" when X = 28 AND Y = 117 else
"100010011101" when X = 29 AND Y = 117 else
"110111011111" when X = 30 AND Y = 117 else
"110111011111" when X = 31 AND Y = 117 else
"110111011111" when X = 32 AND Y = 117 else
"110111011111" when X = 33 AND Y = 117 else
"110111011111" when X = 34 AND Y = 117 else
"110111011111" when X = 35 AND Y = 117 else
"110111011111" when X = 36 AND Y = 117 else
"110111011111" when X = 37 AND Y = 117 else
"110111011111" when X = 38 AND Y = 117 else
"110111011111" when X = 39 AND Y = 117 else
"110111011111" when X = 40 AND Y = 117 else
"110111011111" when X = 41 AND Y = 117 else
"110111011111" when X = 42 AND Y = 117 else
"110111011111" when X = 43 AND Y = 117 else
"110111011111" when X = 44 AND Y = 117 else
"110111011111" when X = 45 AND Y = 117 else
"110111011111" when X = 46 AND Y = 117 else
"110111011111" when X = 47 AND Y = 117 else
"110111011111" when X = 48 AND Y = 117 else
"110111011111" when X = 49 AND Y = 117 else
"110111011111" when X = 50 AND Y = 117 else
"110111011111" when X = 51 AND Y = 117 else
"110111011111" when X = 52 AND Y = 117 else
"110111011111" when X = 53 AND Y = 117 else
"110111011111" when X = 54 AND Y = 117 else
"110111011111" when X = 55 AND Y = 117 else
"110111011111" when X = 56 AND Y = 117 else
"110111011111" when X = 57 AND Y = 117 else
"110111011111" when X = 58 AND Y = 117 else
"110111011111" when X = 59 AND Y = 117 else
"110111011111" when X = 60 AND Y = 117 else
"110111011111" when X = 61 AND Y = 117 else
"110111011111" when X = 62 AND Y = 117 else
"110111011111" when X = 63 AND Y = 117 else
"110111011111" when X = 64 AND Y = 117 else
"110111011111" when X = 65 AND Y = 117 else
"110111011111" when X = 66 AND Y = 117 else
"110111011111" when X = 67 AND Y = 117 else
"110111011111" when X = 68 AND Y = 117 else
"110111011111" when X = 69 AND Y = 117 else
"110111011111" when X = 70 AND Y = 117 else
"110111011111" when X = 71 AND Y = 117 else
"110111011111" when X = 72 AND Y = 117 else
"110111011111" when X = 73 AND Y = 117 else
"110111011111" when X = 74 AND Y = 117 else
"110111011111" when X = 75 AND Y = 117 else
"110111011111" when X = 76 AND Y = 117 else
"110111011111" when X = 77 AND Y = 117 else
"110111011111" when X = 78 AND Y = 117 else
"110111011111" when X = 79 AND Y = 117 else
"110111011111" when X = 80 AND Y = 117 else
"110111011111" when X = 81 AND Y = 117 else
"110111011111" when X = 82 AND Y = 117 else
"110111011111" when X = 83 AND Y = 117 else
"110111011111" when X = 84 AND Y = 117 else
"110111011111" when X = 85 AND Y = 117 else
"110111011111" when X = 86 AND Y = 117 else
"110111011111" when X = 87 AND Y = 117 else
"110111011111" when X = 88 AND Y = 117 else
"110111011111" when X = 89 AND Y = 117 else
"110111011111" when X = 90 AND Y = 117 else
"110111011111" when X = 91 AND Y = 117 else
"110111011111" when X = 92 AND Y = 117 else
"110111011111" when X = 93 AND Y = 117 else
"110111011111" when X = 94 AND Y = 117 else
"110111011111" when X = 95 AND Y = 117 else
"110111011111" when X = 96 AND Y = 117 else
"110111011111" when X = 97 AND Y = 117 else
"110111011111" when X = 98 AND Y = 117 else
"110111011111" when X = 99 AND Y = 117 else
"110111011111" when X = 100 AND Y = 117 else
"110111011111" when X = 101 AND Y = 117 else
"110111011111" when X = 102 AND Y = 117 else
"110111011111" when X = 103 AND Y = 117 else
"110111011111" when X = 104 AND Y = 117 else
"110111011111" when X = 105 AND Y = 117 else
"110111011111" when X = 106 AND Y = 117 else
"110111011111" when X = 107 AND Y = 117 else
"110111011111" when X = 108 AND Y = 117 else
"110111011111" when X = 109 AND Y = 117 else
"110111011111" when X = 110 AND Y = 117 else
"110111011111" when X = 111 AND Y = 117 else
"110111011111" when X = 112 AND Y = 117 else
"110111011111" when X = 113 AND Y = 117 else
"110111011111" when X = 114 AND Y = 117 else
"110111011111" when X = 115 AND Y = 117 else
"110111011111" when X = 116 AND Y = 117 else
"110111011111" when X = 117 AND Y = 117 else
"110111011111" when X = 118 AND Y = 117 else
"110111011111" when X = 119 AND Y = 117 else
"110111011111" when X = 120 AND Y = 117 else
"110111011111" when X = 121 AND Y = 117 else
"110111011111" when X = 122 AND Y = 117 else
"110111011111" when X = 123 AND Y = 117 else
"110111011111" when X = 124 AND Y = 117 else
"110111011111" when X = 125 AND Y = 117 else
"110111011111" when X = 126 AND Y = 117 else
"110111011111" when X = 127 AND Y = 117 else
"110111011111" when X = 128 AND Y = 117 else
"110111011111" when X = 129 AND Y = 117 else
"110111011111" when X = 130 AND Y = 117 else
"110111011111" when X = 131 AND Y = 117 else
"110111011111" when X = 132 AND Y = 117 else
"110111011111" when X = 133 AND Y = 117 else
"110111011111" when X = 134 AND Y = 117 else
"110111011111" when X = 135 AND Y = 117 else
"110111011111" when X = 136 AND Y = 117 else
"110111011111" when X = 137 AND Y = 117 else
"110111011111" when X = 138 AND Y = 117 else
"110111011111" when X = 139 AND Y = 117 else
"110111011111" when X = 140 AND Y = 117 else
"110111011111" when X = 141 AND Y = 117 else
"110111011111" when X = 142 AND Y = 117 else
"110111011111" when X = 143 AND Y = 117 else
"110111011111" when X = 144 AND Y = 117 else
"111111111111" when X = 145 AND Y = 117 else
"111111111111" when X = 146 AND Y = 117 else
"111111111111" when X = 147 AND Y = 117 else
"111111111111" when X = 148 AND Y = 117 else
"111111111111" when X = 149 AND Y = 117 else
"111111111111" when X = 150 AND Y = 117 else
"111111111111" when X = 151 AND Y = 117 else
"111111111111" when X = 152 AND Y = 117 else
"111111111111" when X = 153 AND Y = 117 else
"111111111111" when X = 154 AND Y = 117 else
"111111111111" when X = 155 AND Y = 117 else
"111111111111" when X = 156 AND Y = 117 else
"111111111111" when X = 157 AND Y = 117 else
"111111111111" when X = 158 AND Y = 117 else
"111111111111" when X = 159 AND Y = 117 else
"111111111111" when X = 160 AND Y = 117 else
"111111111111" when X = 161 AND Y = 117 else
"111111111111" when X = 162 AND Y = 117 else
"111111111111" when X = 163 AND Y = 117 else
"111111111111" when X = 164 AND Y = 117 else
"111111111111" when X = 165 AND Y = 117 else
"111111111111" when X = 166 AND Y = 117 else
"111111111111" when X = 167 AND Y = 117 else
"111111111111" when X = 168 AND Y = 117 else
"111111111111" when X = 169 AND Y = 117 else
"111111111111" when X = 170 AND Y = 117 else
"111111111111" when X = 171 AND Y = 117 else
"111111111111" when X = 172 AND Y = 117 else
"111111111111" when X = 173 AND Y = 117 else
"111111111111" when X = 174 AND Y = 117 else
"111111111111" when X = 175 AND Y = 117 else
"111111111111" when X = 176 AND Y = 117 else
"111111111111" when X = 177 AND Y = 117 else
"111111111111" when X = 178 AND Y = 117 else
"111111111111" when X = 179 AND Y = 117 else
"111111111111" when X = 180 AND Y = 117 else
"111111111111" when X = 181 AND Y = 117 else
"111111111111" when X = 182 AND Y = 117 else
"111111111111" when X = 183 AND Y = 117 else
"111111111111" when X = 184 AND Y = 117 else
"111111111111" when X = 185 AND Y = 117 else
"111111111111" when X = 186 AND Y = 117 else
"111111111111" when X = 187 AND Y = 117 else
"111111111111" when X = 188 AND Y = 117 else
"111111111111" when X = 189 AND Y = 117 else
"111111111111" when X = 190 AND Y = 117 else
"111111111111" when X = 191 AND Y = 117 else
"111111111111" when X = 192 AND Y = 117 else
"111111111111" when X = 193 AND Y = 117 else
"111111111111" when X = 194 AND Y = 117 else
"111111111111" when X = 195 AND Y = 117 else
"111111111111" when X = 196 AND Y = 117 else
"111111111111" when X = 197 AND Y = 117 else
"111111111111" when X = 198 AND Y = 117 else
"111111111111" when X = 199 AND Y = 117 else
"111111111111" when X = 200 AND Y = 117 else
"111111111111" when X = 201 AND Y = 117 else
"111111111111" when X = 202 AND Y = 117 else
"111111111111" when X = 203 AND Y = 117 else
"111111111111" when X = 204 AND Y = 117 else
"110111011111" when X = 205 AND Y = 117 else
"110111011111" when X = 206 AND Y = 117 else
"110111011111" when X = 207 AND Y = 117 else
"110111011111" when X = 208 AND Y = 117 else
"110111011111" when X = 209 AND Y = 117 else
"110111011111" when X = 210 AND Y = 117 else
"110111011111" when X = 211 AND Y = 117 else
"110111011111" when X = 212 AND Y = 117 else
"110111011111" when X = 213 AND Y = 117 else
"110111011111" when X = 214 AND Y = 117 else
"110111011111" when X = 215 AND Y = 117 else
"110111011111" when X = 216 AND Y = 117 else
"110111011111" when X = 217 AND Y = 117 else
"110111011111" when X = 218 AND Y = 117 else
"110111011111" when X = 219 AND Y = 117 else
"110111011111" when X = 220 AND Y = 117 else
"110111011111" when X = 221 AND Y = 117 else
"110111011111" when X = 222 AND Y = 117 else
"110111011111" when X = 223 AND Y = 117 else
"110111011111" when X = 224 AND Y = 117 else
"110111011111" when X = 225 AND Y = 117 else
"110111011111" when X = 226 AND Y = 117 else
"110111011111" when X = 227 AND Y = 117 else
"110111011111" when X = 228 AND Y = 117 else
"110111011111" when X = 229 AND Y = 117 else
"110111011111" when X = 230 AND Y = 117 else
"110111011111" when X = 231 AND Y = 117 else
"110111011111" when X = 232 AND Y = 117 else
"110111011111" when X = 233 AND Y = 117 else
"110111011111" when X = 234 AND Y = 117 else
"110111011111" when X = 235 AND Y = 117 else
"110111011111" when X = 236 AND Y = 117 else
"110111011111" when X = 237 AND Y = 117 else
"110111011111" when X = 238 AND Y = 117 else
"110111011111" when X = 239 AND Y = 117 else
"110111011111" when X = 240 AND Y = 117 else
"110111011111" when X = 241 AND Y = 117 else
"110111011111" when X = 242 AND Y = 117 else
"110111011111" when X = 243 AND Y = 117 else
"110111011111" when X = 244 AND Y = 117 else
"110111011111" when X = 245 AND Y = 117 else
"110111011111" when X = 246 AND Y = 117 else
"110111011111" when X = 247 AND Y = 117 else
"110111011111" when X = 248 AND Y = 117 else
"110111011111" when X = 249 AND Y = 117 else
"110111011111" when X = 250 AND Y = 117 else
"110111011111" when X = 251 AND Y = 117 else
"110111011111" when X = 252 AND Y = 117 else
"110111011111" when X = 253 AND Y = 117 else
"110111011111" when X = 254 AND Y = 117 else
"110111011111" when X = 255 AND Y = 117 else
"110111011111" when X = 256 AND Y = 117 else
"110111011111" when X = 257 AND Y = 117 else
"110111011111" when X = 258 AND Y = 117 else
"110111011111" when X = 259 AND Y = 117 else
"110111011111" when X = 260 AND Y = 117 else
"110111011111" when X = 261 AND Y = 117 else
"110111011111" when X = 262 AND Y = 117 else
"110111011111" when X = 263 AND Y = 117 else
"110111011111" when X = 264 AND Y = 117 else
"110111011111" when X = 265 AND Y = 117 else
"110111011111" when X = 266 AND Y = 117 else
"110111011111" when X = 267 AND Y = 117 else
"110111011111" when X = 268 AND Y = 117 else
"110111011111" when X = 269 AND Y = 117 else
"110111011111" when X = 270 AND Y = 117 else
"110111011111" when X = 271 AND Y = 117 else
"110111011111" when X = 272 AND Y = 117 else
"110111011111" when X = 273 AND Y = 117 else
"110111011111" when X = 274 AND Y = 117 else
"110111011111" when X = 275 AND Y = 117 else
"110111011111" when X = 276 AND Y = 117 else
"110111011111" when X = 277 AND Y = 117 else
"110111011111" when X = 278 AND Y = 117 else
"110111011111" when X = 279 AND Y = 117 else
"111111111111" when X = 280 AND Y = 117 else
"111111111111" when X = 281 AND Y = 117 else
"111111111111" when X = 282 AND Y = 117 else
"111111111111" when X = 283 AND Y = 117 else
"111111111111" when X = 284 AND Y = 117 else
"111111111111" when X = 285 AND Y = 117 else
"111111111111" when X = 286 AND Y = 117 else
"111111111111" when X = 287 AND Y = 117 else
"111111111111" when X = 288 AND Y = 117 else
"111111111111" when X = 289 AND Y = 117 else
"111111111111" when X = 290 AND Y = 117 else
"111111111111" when X = 291 AND Y = 117 else
"111111111111" when X = 292 AND Y = 117 else
"111111111111" when X = 293 AND Y = 117 else
"111111111111" when X = 294 AND Y = 117 else
"111111111111" when X = 295 AND Y = 117 else
"111111111111" when X = 296 AND Y = 117 else
"111111111111" when X = 297 AND Y = 117 else
"111111111111" when X = 298 AND Y = 117 else
"111111111111" when X = 299 AND Y = 117 else
"110111011111" when X = 300 AND Y = 117 else
"110111011111" when X = 301 AND Y = 117 else
"110111011111" when X = 302 AND Y = 117 else
"110111011111" when X = 303 AND Y = 117 else
"110111011111" when X = 304 AND Y = 117 else
"110111011111" when X = 305 AND Y = 117 else
"110111011111" when X = 306 AND Y = 117 else
"110111011111" when X = 307 AND Y = 117 else
"110111011111" when X = 308 AND Y = 117 else
"110111011111" when X = 309 AND Y = 117 else
"110111011111" when X = 310 AND Y = 117 else
"110111011111" when X = 311 AND Y = 117 else
"110111011111" when X = 312 AND Y = 117 else
"110111011111" when X = 313 AND Y = 117 else
"110111011111" when X = 314 AND Y = 117 else
"110111011111" when X = 315 AND Y = 117 else
"110111011111" when X = 316 AND Y = 117 else
"110111011111" when X = 317 AND Y = 117 else
"110111011111" when X = 318 AND Y = 117 else
"110111011111" when X = 319 AND Y = 117 else
"110111011111" when X = 320 AND Y = 117 else
"110111011111" when X = 321 AND Y = 117 else
"110111011111" when X = 322 AND Y = 117 else
"110111011111" when X = 323 AND Y = 117 else
"110111011111" when X = 324 AND Y = 117 else
"100010011101" when X = 0 AND Y = 118 else
"100010011101" when X = 1 AND Y = 118 else
"100010011101" when X = 2 AND Y = 118 else
"100010011101" when X = 3 AND Y = 118 else
"100010011101" when X = 4 AND Y = 118 else
"100010011101" when X = 5 AND Y = 118 else
"100010011101" when X = 6 AND Y = 118 else
"100010011101" when X = 7 AND Y = 118 else
"100010011101" when X = 8 AND Y = 118 else
"100010011101" when X = 9 AND Y = 118 else
"100010011101" when X = 10 AND Y = 118 else
"100010011101" when X = 11 AND Y = 118 else
"100010011101" when X = 12 AND Y = 118 else
"100010011101" when X = 13 AND Y = 118 else
"100010011101" when X = 14 AND Y = 118 else
"100010011101" when X = 15 AND Y = 118 else
"100010011101" when X = 16 AND Y = 118 else
"100010011101" when X = 17 AND Y = 118 else
"100010011101" when X = 18 AND Y = 118 else
"100010011101" when X = 19 AND Y = 118 else
"100010011101" when X = 20 AND Y = 118 else
"100010011101" when X = 21 AND Y = 118 else
"100010011101" when X = 22 AND Y = 118 else
"100010011101" when X = 23 AND Y = 118 else
"100010011101" when X = 24 AND Y = 118 else
"100010011101" when X = 25 AND Y = 118 else
"100010011101" when X = 26 AND Y = 118 else
"100010011101" when X = 27 AND Y = 118 else
"100010011101" when X = 28 AND Y = 118 else
"100010011101" when X = 29 AND Y = 118 else
"110111011111" when X = 30 AND Y = 118 else
"110111011111" when X = 31 AND Y = 118 else
"110111011111" when X = 32 AND Y = 118 else
"110111011111" when X = 33 AND Y = 118 else
"110111011111" when X = 34 AND Y = 118 else
"110111011111" when X = 35 AND Y = 118 else
"110111011111" when X = 36 AND Y = 118 else
"110111011111" when X = 37 AND Y = 118 else
"110111011111" when X = 38 AND Y = 118 else
"110111011111" when X = 39 AND Y = 118 else
"110111011111" when X = 40 AND Y = 118 else
"110111011111" when X = 41 AND Y = 118 else
"110111011111" when X = 42 AND Y = 118 else
"110111011111" when X = 43 AND Y = 118 else
"110111011111" when X = 44 AND Y = 118 else
"110111011111" when X = 45 AND Y = 118 else
"110111011111" when X = 46 AND Y = 118 else
"110111011111" when X = 47 AND Y = 118 else
"110111011111" when X = 48 AND Y = 118 else
"110111011111" when X = 49 AND Y = 118 else
"110111011111" when X = 50 AND Y = 118 else
"110111011111" when X = 51 AND Y = 118 else
"110111011111" when X = 52 AND Y = 118 else
"110111011111" when X = 53 AND Y = 118 else
"110111011111" when X = 54 AND Y = 118 else
"110111011111" when X = 55 AND Y = 118 else
"110111011111" when X = 56 AND Y = 118 else
"110111011111" when X = 57 AND Y = 118 else
"110111011111" when X = 58 AND Y = 118 else
"110111011111" when X = 59 AND Y = 118 else
"110111011111" when X = 60 AND Y = 118 else
"110111011111" when X = 61 AND Y = 118 else
"110111011111" when X = 62 AND Y = 118 else
"110111011111" when X = 63 AND Y = 118 else
"110111011111" when X = 64 AND Y = 118 else
"110111011111" when X = 65 AND Y = 118 else
"110111011111" when X = 66 AND Y = 118 else
"110111011111" when X = 67 AND Y = 118 else
"110111011111" when X = 68 AND Y = 118 else
"110111011111" when X = 69 AND Y = 118 else
"110111011111" when X = 70 AND Y = 118 else
"110111011111" when X = 71 AND Y = 118 else
"110111011111" when X = 72 AND Y = 118 else
"110111011111" when X = 73 AND Y = 118 else
"110111011111" when X = 74 AND Y = 118 else
"110111011111" when X = 75 AND Y = 118 else
"110111011111" when X = 76 AND Y = 118 else
"110111011111" when X = 77 AND Y = 118 else
"110111011111" when X = 78 AND Y = 118 else
"110111011111" when X = 79 AND Y = 118 else
"110111011111" when X = 80 AND Y = 118 else
"110111011111" when X = 81 AND Y = 118 else
"110111011111" when X = 82 AND Y = 118 else
"110111011111" when X = 83 AND Y = 118 else
"110111011111" when X = 84 AND Y = 118 else
"110111011111" when X = 85 AND Y = 118 else
"110111011111" when X = 86 AND Y = 118 else
"110111011111" when X = 87 AND Y = 118 else
"110111011111" when X = 88 AND Y = 118 else
"110111011111" when X = 89 AND Y = 118 else
"110111011111" when X = 90 AND Y = 118 else
"110111011111" when X = 91 AND Y = 118 else
"110111011111" when X = 92 AND Y = 118 else
"110111011111" when X = 93 AND Y = 118 else
"110111011111" when X = 94 AND Y = 118 else
"110111011111" when X = 95 AND Y = 118 else
"110111011111" when X = 96 AND Y = 118 else
"110111011111" when X = 97 AND Y = 118 else
"110111011111" when X = 98 AND Y = 118 else
"110111011111" when X = 99 AND Y = 118 else
"110111011111" when X = 100 AND Y = 118 else
"110111011111" when X = 101 AND Y = 118 else
"110111011111" when X = 102 AND Y = 118 else
"110111011111" when X = 103 AND Y = 118 else
"110111011111" when X = 104 AND Y = 118 else
"110111011111" when X = 105 AND Y = 118 else
"110111011111" when X = 106 AND Y = 118 else
"110111011111" when X = 107 AND Y = 118 else
"110111011111" when X = 108 AND Y = 118 else
"110111011111" when X = 109 AND Y = 118 else
"110111011111" when X = 110 AND Y = 118 else
"110111011111" when X = 111 AND Y = 118 else
"110111011111" when X = 112 AND Y = 118 else
"110111011111" when X = 113 AND Y = 118 else
"110111011111" when X = 114 AND Y = 118 else
"110111011111" when X = 115 AND Y = 118 else
"110111011111" when X = 116 AND Y = 118 else
"110111011111" when X = 117 AND Y = 118 else
"110111011111" when X = 118 AND Y = 118 else
"110111011111" when X = 119 AND Y = 118 else
"110111011111" when X = 120 AND Y = 118 else
"110111011111" when X = 121 AND Y = 118 else
"110111011111" when X = 122 AND Y = 118 else
"110111011111" when X = 123 AND Y = 118 else
"110111011111" when X = 124 AND Y = 118 else
"110111011111" when X = 125 AND Y = 118 else
"110111011111" when X = 126 AND Y = 118 else
"110111011111" when X = 127 AND Y = 118 else
"110111011111" when X = 128 AND Y = 118 else
"110111011111" when X = 129 AND Y = 118 else
"110111011111" when X = 130 AND Y = 118 else
"110111011111" when X = 131 AND Y = 118 else
"110111011111" when X = 132 AND Y = 118 else
"110111011111" when X = 133 AND Y = 118 else
"110111011111" when X = 134 AND Y = 118 else
"110111011111" when X = 135 AND Y = 118 else
"110111011111" when X = 136 AND Y = 118 else
"110111011111" when X = 137 AND Y = 118 else
"110111011111" when X = 138 AND Y = 118 else
"110111011111" when X = 139 AND Y = 118 else
"110111011111" when X = 140 AND Y = 118 else
"110111011111" when X = 141 AND Y = 118 else
"110111011111" when X = 142 AND Y = 118 else
"110111011111" when X = 143 AND Y = 118 else
"110111011111" when X = 144 AND Y = 118 else
"111111111111" when X = 145 AND Y = 118 else
"111111111111" when X = 146 AND Y = 118 else
"111111111111" when X = 147 AND Y = 118 else
"111111111111" when X = 148 AND Y = 118 else
"111111111111" when X = 149 AND Y = 118 else
"111111111111" when X = 150 AND Y = 118 else
"111111111111" when X = 151 AND Y = 118 else
"111111111111" when X = 152 AND Y = 118 else
"111111111111" when X = 153 AND Y = 118 else
"111111111111" when X = 154 AND Y = 118 else
"111111111111" when X = 155 AND Y = 118 else
"111111111111" when X = 156 AND Y = 118 else
"111111111111" when X = 157 AND Y = 118 else
"111111111111" when X = 158 AND Y = 118 else
"111111111111" when X = 159 AND Y = 118 else
"111111111111" when X = 160 AND Y = 118 else
"111111111111" when X = 161 AND Y = 118 else
"111111111111" when X = 162 AND Y = 118 else
"111111111111" when X = 163 AND Y = 118 else
"111111111111" when X = 164 AND Y = 118 else
"111111111111" when X = 165 AND Y = 118 else
"111111111111" when X = 166 AND Y = 118 else
"111111111111" when X = 167 AND Y = 118 else
"111111111111" when X = 168 AND Y = 118 else
"111111111111" when X = 169 AND Y = 118 else
"111111111111" when X = 170 AND Y = 118 else
"111111111111" when X = 171 AND Y = 118 else
"111111111111" when X = 172 AND Y = 118 else
"111111111111" when X = 173 AND Y = 118 else
"111111111111" when X = 174 AND Y = 118 else
"111111111111" when X = 175 AND Y = 118 else
"111111111111" when X = 176 AND Y = 118 else
"111111111111" when X = 177 AND Y = 118 else
"111111111111" when X = 178 AND Y = 118 else
"111111111111" when X = 179 AND Y = 118 else
"111111111111" when X = 180 AND Y = 118 else
"111111111111" when X = 181 AND Y = 118 else
"111111111111" when X = 182 AND Y = 118 else
"111111111111" when X = 183 AND Y = 118 else
"111111111111" when X = 184 AND Y = 118 else
"111111111111" when X = 185 AND Y = 118 else
"111111111111" when X = 186 AND Y = 118 else
"111111111111" when X = 187 AND Y = 118 else
"111111111111" when X = 188 AND Y = 118 else
"111111111111" when X = 189 AND Y = 118 else
"111111111111" when X = 190 AND Y = 118 else
"111111111111" when X = 191 AND Y = 118 else
"111111111111" when X = 192 AND Y = 118 else
"111111111111" when X = 193 AND Y = 118 else
"111111111111" when X = 194 AND Y = 118 else
"111111111111" when X = 195 AND Y = 118 else
"111111111111" when X = 196 AND Y = 118 else
"111111111111" when X = 197 AND Y = 118 else
"111111111111" when X = 198 AND Y = 118 else
"111111111111" when X = 199 AND Y = 118 else
"111111111111" when X = 200 AND Y = 118 else
"111111111111" when X = 201 AND Y = 118 else
"111111111111" when X = 202 AND Y = 118 else
"111111111111" when X = 203 AND Y = 118 else
"111111111111" when X = 204 AND Y = 118 else
"110111011111" when X = 205 AND Y = 118 else
"110111011111" when X = 206 AND Y = 118 else
"110111011111" when X = 207 AND Y = 118 else
"110111011111" when X = 208 AND Y = 118 else
"110111011111" when X = 209 AND Y = 118 else
"110111011111" when X = 210 AND Y = 118 else
"110111011111" when X = 211 AND Y = 118 else
"110111011111" when X = 212 AND Y = 118 else
"110111011111" when X = 213 AND Y = 118 else
"110111011111" when X = 214 AND Y = 118 else
"110111011111" when X = 215 AND Y = 118 else
"110111011111" when X = 216 AND Y = 118 else
"110111011111" when X = 217 AND Y = 118 else
"110111011111" when X = 218 AND Y = 118 else
"110111011111" when X = 219 AND Y = 118 else
"110111011111" when X = 220 AND Y = 118 else
"110111011111" when X = 221 AND Y = 118 else
"110111011111" when X = 222 AND Y = 118 else
"110111011111" when X = 223 AND Y = 118 else
"110111011111" when X = 224 AND Y = 118 else
"110111011111" when X = 225 AND Y = 118 else
"110111011111" when X = 226 AND Y = 118 else
"110111011111" when X = 227 AND Y = 118 else
"110111011111" when X = 228 AND Y = 118 else
"110111011111" when X = 229 AND Y = 118 else
"110111011111" when X = 230 AND Y = 118 else
"110111011111" when X = 231 AND Y = 118 else
"110111011111" when X = 232 AND Y = 118 else
"110111011111" when X = 233 AND Y = 118 else
"110111011111" when X = 234 AND Y = 118 else
"110111011111" when X = 235 AND Y = 118 else
"110111011111" when X = 236 AND Y = 118 else
"110111011111" when X = 237 AND Y = 118 else
"110111011111" when X = 238 AND Y = 118 else
"110111011111" when X = 239 AND Y = 118 else
"110111011111" when X = 240 AND Y = 118 else
"110111011111" when X = 241 AND Y = 118 else
"110111011111" when X = 242 AND Y = 118 else
"110111011111" when X = 243 AND Y = 118 else
"110111011111" when X = 244 AND Y = 118 else
"110111011111" when X = 245 AND Y = 118 else
"110111011111" when X = 246 AND Y = 118 else
"110111011111" when X = 247 AND Y = 118 else
"110111011111" when X = 248 AND Y = 118 else
"110111011111" when X = 249 AND Y = 118 else
"110111011111" when X = 250 AND Y = 118 else
"110111011111" when X = 251 AND Y = 118 else
"110111011111" when X = 252 AND Y = 118 else
"110111011111" when X = 253 AND Y = 118 else
"110111011111" when X = 254 AND Y = 118 else
"110111011111" when X = 255 AND Y = 118 else
"110111011111" when X = 256 AND Y = 118 else
"110111011111" when X = 257 AND Y = 118 else
"110111011111" when X = 258 AND Y = 118 else
"110111011111" when X = 259 AND Y = 118 else
"110111011111" when X = 260 AND Y = 118 else
"110111011111" when X = 261 AND Y = 118 else
"110111011111" when X = 262 AND Y = 118 else
"110111011111" when X = 263 AND Y = 118 else
"110111011111" when X = 264 AND Y = 118 else
"110111011111" when X = 265 AND Y = 118 else
"110111011111" when X = 266 AND Y = 118 else
"110111011111" when X = 267 AND Y = 118 else
"110111011111" when X = 268 AND Y = 118 else
"110111011111" when X = 269 AND Y = 118 else
"110111011111" when X = 270 AND Y = 118 else
"110111011111" when X = 271 AND Y = 118 else
"110111011111" when X = 272 AND Y = 118 else
"110111011111" when X = 273 AND Y = 118 else
"110111011111" when X = 274 AND Y = 118 else
"110111011111" when X = 275 AND Y = 118 else
"110111011111" when X = 276 AND Y = 118 else
"110111011111" when X = 277 AND Y = 118 else
"110111011111" when X = 278 AND Y = 118 else
"110111011111" when X = 279 AND Y = 118 else
"111111111111" when X = 280 AND Y = 118 else
"111111111111" when X = 281 AND Y = 118 else
"111111111111" when X = 282 AND Y = 118 else
"111111111111" when X = 283 AND Y = 118 else
"111111111111" when X = 284 AND Y = 118 else
"111111111111" when X = 285 AND Y = 118 else
"111111111111" when X = 286 AND Y = 118 else
"111111111111" when X = 287 AND Y = 118 else
"111111111111" when X = 288 AND Y = 118 else
"111111111111" when X = 289 AND Y = 118 else
"111111111111" when X = 290 AND Y = 118 else
"111111111111" when X = 291 AND Y = 118 else
"111111111111" when X = 292 AND Y = 118 else
"111111111111" when X = 293 AND Y = 118 else
"111111111111" when X = 294 AND Y = 118 else
"111111111111" when X = 295 AND Y = 118 else
"111111111111" when X = 296 AND Y = 118 else
"111111111111" when X = 297 AND Y = 118 else
"111111111111" when X = 298 AND Y = 118 else
"111111111111" when X = 299 AND Y = 118 else
"110111011111" when X = 300 AND Y = 118 else
"110111011111" when X = 301 AND Y = 118 else
"110111011111" when X = 302 AND Y = 118 else
"110111011111" when X = 303 AND Y = 118 else
"110111011111" when X = 304 AND Y = 118 else
"110111011111" when X = 305 AND Y = 118 else
"110111011111" when X = 306 AND Y = 118 else
"110111011111" when X = 307 AND Y = 118 else
"110111011111" when X = 308 AND Y = 118 else
"110111011111" when X = 309 AND Y = 118 else
"110111011111" when X = 310 AND Y = 118 else
"110111011111" when X = 311 AND Y = 118 else
"110111011111" when X = 312 AND Y = 118 else
"110111011111" when X = 313 AND Y = 118 else
"110111011111" when X = 314 AND Y = 118 else
"110111011111" when X = 315 AND Y = 118 else
"110111011111" when X = 316 AND Y = 118 else
"110111011111" when X = 317 AND Y = 118 else
"110111011111" when X = 318 AND Y = 118 else
"110111011111" when X = 319 AND Y = 118 else
"110111011111" when X = 320 AND Y = 118 else
"110111011111" when X = 321 AND Y = 118 else
"110111011111" when X = 322 AND Y = 118 else
"110111011111" when X = 323 AND Y = 118 else
"110111011111" when X = 324 AND Y = 118 else
"100010011101" when X = 0 AND Y = 119 else
"100010011101" when X = 1 AND Y = 119 else
"100010011101" when X = 2 AND Y = 119 else
"100010011101" when X = 3 AND Y = 119 else
"100010011101" when X = 4 AND Y = 119 else
"100010011101" when X = 5 AND Y = 119 else
"100010011101" when X = 6 AND Y = 119 else
"100010011101" when X = 7 AND Y = 119 else
"100010011101" when X = 8 AND Y = 119 else
"100010011101" when X = 9 AND Y = 119 else
"100010011101" when X = 10 AND Y = 119 else
"100010011101" when X = 11 AND Y = 119 else
"100010011101" when X = 12 AND Y = 119 else
"100010011101" when X = 13 AND Y = 119 else
"100010011101" when X = 14 AND Y = 119 else
"100010011101" when X = 15 AND Y = 119 else
"100010011101" when X = 16 AND Y = 119 else
"100010011101" when X = 17 AND Y = 119 else
"100010011101" when X = 18 AND Y = 119 else
"100010011101" when X = 19 AND Y = 119 else
"100010011101" when X = 20 AND Y = 119 else
"100010011101" when X = 21 AND Y = 119 else
"100010011101" when X = 22 AND Y = 119 else
"100010011101" when X = 23 AND Y = 119 else
"100010011101" when X = 24 AND Y = 119 else
"100010011101" when X = 25 AND Y = 119 else
"100010011101" when X = 26 AND Y = 119 else
"100010011101" when X = 27 AND Y = 119 else
"100010011101" when X = 28 AND Y = 119 else
"100010011101" when X = 29 AND Y = 119 else
"110111011111" when X = 30 AND Y = 119 else
"110111011111" when X = 31 AND Y = 119 else
"110111011111" when X = 32 AND Y = 119 else
"110111011111" when X = 33 AND Y = 119 else
"110111011111" when X = 34 AND Y = 119 else
"110111011111" when X = 35 AND Y = 119 else
"110111011111" when X = 36 AND Y = 119 else
"110111011111" when X = 37 AND Y = 119 else
"110111011111" when X = 38 AND Y = 119 else
"110111011111" when X = 39 AND Y = 119 else
"110111011111" when X = 40 AND Y = 119 else
"110111011111" when X = 41 AND Y = 119 else
"110111011111" when X = 42 AND Y = 119 else
"110111011111" when X = 43 AND Y = 119 else
"110111011111" when X = 44 AND Y = 119 else
"110111011111" when X = 45 AND Y = 119 else
"110111011111" when X = 46 AND Y = 119 else
"110111011111" when X = 47 AND Y = 119 else
"110111011111" when X = 48 AND Y = 119 else
"110111011111" when X = 49 AND Y = 119 else
"110111011111" when X = 50 AND Y = 119 else
"110111011111" when X = 51 AND Y = 119 else
"110111011111" when X = 52 AND Y = 119 else
"110111011111" when X = 53 AND Y = 119 else
"110111011111" when X = 54 AND Y = 119 else
"110111011111" when X = 55 AND Y = 119 else
"110111011111" when X = 56 AND Y = 119 else
"110111011111" when X = 57 AND Y = 119 else
"110111011111" when X = 58 AND Y = 119 else
"110111011111" when X = 59 AND Y = 119 else
"110111011111" when X = 60 AND Y = 119 else
"110111011111" when X = 61 AND Y = 119 else
"110111011111" when X = 62 AND Y = 119 else
"110111011111" when X = 63 AND Y = 119 else
"110111011111" when X = 64 AND Y = 119 else
"110111011111" when X = 65 AND Y = 119 else
"110111011111" when X = 66 AND Y = 119 else
"110111011111" when X = 67 AND Y = 119 else
"110111011111" when X = 68 AND Y = 119 else
"110111011111" when X = 69 AND Y = 119 else
"110111011111" when X = 70 AND Y = 119 else
"110111011111" when X = 71 AND Y = 119 else
"110111011111" when X = 72 AND Y = 119 else
"110111011111" when X = 73 AND Y = 119 else
"110111011111" when X = 74 AND Y = 119 else
"110111011111" when X = 75 AND Y = 119 else
"110111011111" when X = 76 AND Y = 119 else
"110111011111" when X = 77 AND Y = 119 else
"110111011111" when X = 78 AND Y = 119 else
"110111011111" when X = 79 AND Y = 119 else
"110111011111" when X = 80 AND Y = 119 else
"110111011111" when X = 81 AND Y = 119 else
"110111011111" when X = 82 AND Y = 119 else
"110111011111" when X = 83 AND Y = 119 else
"110111011111" when X = 84 AND Y = 119 else
"110111011111" when X = 85 AND Y = 119 else
"110111011111" when X = 86 AND Y = 119 else
"110111011111" when X = 87 AND Y = 119 else
"110111011111" when X = 88 AND Y = 119 else
"110111011111" when X = 89 AND Y = 119 else
"110111011111" when X = 90 AND Y = 119 else
"110111011111" when X = 91 AND Y = 119 else
"110111011111" when X = 92 AND Y = 119 else
"110111011111" when X = 93 AND Y = 119 else
"110111011111" when X = 94 AND Y = 119 else
"110111011111" when X = 95 AND Y = 119 else
"110111011111" when X = 96 AND Y = 119 else
"110111011111" when X = 97 AND Y = 119 else
"110111011111" when X = 98 AND Y = 119 else
"110111011111" when X = 99 AND Y = 119 else
"110111011111" when X = 100 AND Y = 119 else
"110111011111" when X = 101 AND Y = 119 else
"110111011111" when X = 102 AND Y = 119 else
"110111011111" when X = 103 AND Y = 119 else
"110111011111" when X = 104 AND Y = 119 else
"110111011111" when X = 105 AND Y = 119 else
"110111011111" when X = 106 AND Y = 119 else
"110111011111" when X = 107 AND Y = 119 else
"110111011111" when X = 108 AND Y = 119 else
"110111011111" when X = 109 AND Y = 119 else
"110111011111" when X = 110 AND Y = 119 else
"110111011111" when X = 111 AND Y = 119 else
"110111011111" when X = 112 AND Y = 119 else
"110111011111" when X = 113 AND Y = 119 else
"110111011111" when X = 114 AND Y = 119 else
"110111011111" when X = 115 AND Y = 119 else
"110111011111" when X = 116 AND Y = 119 else
"110111011111" when X = 117 AND Y = 119 else
"110111011111" when X = 118 AND Y = 119 else
"110111011111" when X = 119 AND Y = 119 else
"110111011111" when X = 120 AND Y = 119 else
"110111011111" when X = 121 AND Y = 119 else
"110111011111" when X = 122 AND Y = 119 else
"110111011111" when X = 123 AND Y = 119 else
"110111011111" when X = 124 AND Y = 119 else
"110111011111" when X = 125 AND Y = 119 else
"110111011111" when X = 126 AND Y = 119 else
"110111011111" when X = 127 AND Y = 119 else
"110111011111" when X = 128 AND Y = 119 else
"110111011111" when X = 129 AND Y = 119 else
"110111011111" when X = 130 AND Y = 119 else
"110111011111" when X = 131 AND Y = 119 else
"110111011111" when X = 132 AND Y = 119 else
"110111011111" when X = 133 AND Y = 119 else
"110111011111" when X = 134 AND Y = 119 else
"110111011111" when X = 135 AND Y = 119 else
"110111011111" when X = 136 AND Y = 119 else
"110111011111" when X = 137 AND Y = 119 else
"110111011111" when X = 138 AND Y = 119 else
"110111011111" when X = 139 AND Y = 119 else
"110111011111" when X = 140 AND Y = 119 else
"110111011111" when X = 141 AND Y = 119 else
"110111011111" when X = 142 AND Y = 119 else
"110111011111" when X = 143 AND Y = 119 else
"110111011111" when X = 144 AND Y = 119 else
"111111111111" when X = 145 AND Y = 119 else
"111111111111" when X = 146 AND Y = 119 else
"111111111111" when X = 147 AND Y = 119 else
"111111111111" when X = 148 AND Y = 119 else
"111111111111" when X = 149 AND Y = 119 else
"111111111111" when X = 150 AND Y = 119 else
"111111111111" when X = 151 AND Y = 119 else
"111111111111" when X = 152 AND Y = 119 else
"111111111111" when X = 153 AND Y = 119 else
"111111111111" when X = 154 AND Y = 119 else
"111111111111" when X = 155 AND Y = 119 else
"111111111111" when X = 156 AND Y = 119 else
"111111111111" when X = 157 AND Y = 119 else
"111111111111" when X = 158 AND Y = 119 else
"111111111111" when X = 159 AND Y = 119 else
"111111111111" when X = 160 AND Y = 119 else
"111111111111" when X = 161 AND Y = 119 else
"111111111111" when X = 162 AND Y = 119 else
"111111111111" when X = 163 AND Y = 119 else
"111111111111" when X = 164 AND Y = 119 else
"111111111111" when X = 165 AND Y = 119 else
"111111111111" when X = 166 AND Y = 119 else
"111111111111" when X = 167 AND Y = 119 else
"111111111111" when X = 168 AND Y = 119 else
"111111111111" when X = 169 AND Y = 119 else
"111111111111" when X = 170 AND Y = 119 else
"111111111111" when X = 171 AND Y = 119 else
"111111111111" when X = 172 AND Y = 119 else
"111111111111" when X = 173 AND Y = 119 else
"111111111111" when X = 174 AND Y = 119 else
"111111111111" when X = 175 AND Y = 119 else
"111111111111" when X = 176 AND Y = 119 else
"111111111111" when X = 177 AND Y = 119 else
"111111111111" when X = 178 AND Y = 119 else
"111111111111" when X = 179 AND Y = 119 else
"111111111111" when X = 180 AND Y = 119 else
"111111111111" when X = 181 AND Y = 119 else
"111111111111" when X = 182 AND Y = 119 else
"111111111111" when X = 183 AND Y = 119 else
"111111111111" when X = 184 AND Y = 119 else
"111111111111" when X = 185 AND Y = 119 else
"111111111111" when X = 186 AND Y = 119 else
"111111111111" when X = 187 AND Y = 119 else
"111111111111" when X = 188 AND Y = 119 else
"111111111111" when X = 189 AND Y = 119 else
"111111111111" when X = 190 AND Y = 119 else
"111111111111" when X = 191 AND Y = 119 else
"111111111111" when X = 192 AND Y = 119 else
"111111111111" when X = 193 AND Y = 119 else
"111111111111" when X = 194 AND Y = 119 else
"111111111111" when X = 195 AND Y = 119 else
"111111111111" when X = 196 AND Y = 119 else
"111111111111" when X = 197 AND Y = 119 else
"111111111111" when X = 198 AND Y = 119 else
"111111111111" when X = 199 AND Y = 119 else
"111111111111" when X = 200 AND Y = 119 else
"111111111111" when X = 201 AND Y = 119 else
"111111111111" when X = 202 AND Y = 119 else
"111111111111" when X = 203 AND Y = 119 else
"111111111111" when X = 204 AND Y = 119 else
"110111011111" when X = 205 AND Y = 119 else
"110111011111" when X = 206 AND Y = 119 else
"110111011111" when X = 207 AND Y = 119 else
"110111011111" when X = 208 AND Y = 119 else
"110111011111" when X = 209 AND Y = 119 else
"110111011111" when X = 210 AND Y = 119 else
"110111011111" when X = 211 AND Y = 119 else
"110111011111" when X = 212 AND Y = 119 else
"110111011111" when X = 213 AND Y = 119 else
"110111011111" when X = 214 AND Y = 119 else
"110111011111" when X = 215 AND Y = 119 else
"110111011111" when X = 216 AND Y = 119 else
"110111011111" when X = 217 AND Y = 119 else
"110111011111" when X = 218 AND Y = 119 else
"110111011111" when X = 219 AND Y = 119 else
"110111011111" when X = 220 AND Y = 119 else
"110111011111" when X = 221 AND Y = 119 else
"110111011111" when X = 222 AND Y = 119 else
"110111011111" when X = 223 AND Y = 119 else
"110111011111" when X = 224 AND Y = 119 else
"110111011111" when X = 225 AND Y = 119 else
"110111011111" when X = 226 AND Y = 119 else
"110111011111" when X = 227 AND Y = 119 else
"110111011111" when X = 228 AND Y = 119 else
"110111011111" when X = 229 AND Y = 119 else
"110111011111" when X = 230 AND Y = 119 else
"110111011111" when X = 231 AND Y = 119 else
"110111011111" when X = 232 AND Y = 119 else
"110111011111" when X = 233 AND Y = 119 else
"110111011111" when X = 234 AND Y = 119 else
"110111011111" when X = 235 AND Y = 119 else
"110111011111" when X = 236 AND Y = 119 else
"110111011111" when X = 237 AND Y = 119 else
"110111011111" when X = 238 AND Y = 119 else
"110111011111" when X = 239 AND Y = 119 else
"110111011111" when X = 240 AND Y = 119 else
"110111011111" when X = 241 AND Y = 119 else
"110111011111" when X = 242 AND Y = 119 else
"110111011111" when X = 243 AND Y = 119 else
"110111011111" when X = 244 AND Y = 119 else
"110111011111" when X = 245 AND Y = 119 else
"110111011111" when X = 246 AND Y = 119 else
"110111011111" when X = 247 AND Y = 119 else
"110111011111" when X = 248 AND Y = 119 else
"110111011111" when X = 249 AND Y = 119 else
"110111011111" when X = 250 AND Y = 119 else
"110111011111" when X = 251 AND Y = 119 else
"110111011111" when X = 252 AND Y = 119 else
"110111011111" when X = 253 AND Y = 119 else
"110111011111" when X = 254 AND Y = 119 else
"110111011111" when X = 255 AND Y = 119 else
"110111011111" when X = 256 AND Y = 119 else
"110111011111" when X = 257 AND Y = 119 else
"110111011111" when X = 258 AND Y = 119 else
"110111011111" when X = 259 AND Y = 119 else
"110111011111" when X = 260 AND Y = 119 else
"110111011111" when X = 261 AND Y = 119 else
"110111011111" when X = 262 AND Y = 119 else
"110111011111" when X = 263 AND Y = 119 else
"110111011111" when X = 264 AND Y = 119 else
"110111011111" when X = 265 AND Y = 119 else
"110111011111" when X = 266 AND Y = 119 else
"110111011111" when X = 267 AND Y = 119 else
"110111011111" when X = 268 AND Y = 119 else
"110111011111" when X = 269 AND Y = 119 else
"110111011111" when X = 270 AND Y = 119 else
"110111011111" when X = 271 AND Y = 119 else
"110111011111" when X = 272 AND Y = 119 else
"110111011111" when X = 273 AND Y = 119 else
"110111011111" when X = 274 AND Y = 119 else
"110111011111" when X = 275 AND Y = 119 else
"110111011111" when X = 276 AND Y = 119 else
"110111011111" when X = 277 AND Y = 119 else
"110111011111" when X = 278 AND Y = 119 else
"110111011111" when X = 279 AND Y = 119 else
"111111111111" when X = 280 AND Y = 119 else
"111111111111" when X = 281 AND Y = 119 else
"111111111111" when X = 282 AND Y = 119 else
"111111111111" when X = 283 AND Y = 119 else
"111111111111" when X = 284 AND Y = 119 else
"111111111111" when X = 285 AND Y = 119 else
"111111111111" when X = 286 AND Y = 119 else
"111111111111" when X = 287 AND Y = 119 else
"111111111111" when X = 288 AND Y = 119 else
"111111111111" when X = 289 AND Y = 119 else
"111111111111" when X = 290 AND Y = 119 else
"111111111111" when X = 291 AND Y = 119 else
"111111111111" when X = 292 AND Y = 119 else
"111111111111" when X = 293 AND Y = 119 else
"111111111111" when X = 294 AND Y = 119 else
"111111111111" when X = 295 AND Y = 119 else
"111111111111" when X = 296 AND Y = 119 else
"111111111111" when X = 297 AND Y = 119 else
"111111111111" when X = 298 AND Y = 119 else
"111111111111" when X = 299 AND Y = 119 else
"110111011111" when X = 300 AND Y = 119 else
"110111011111" when X = 301 AND Y = 119 else
"110111011111" when X = 302 AND Y = 119 else
"110111011111" when X = 303 AND Y = 119 else
"110111011111" when X = 304 AND Y = 119 else
"110111011111" when X = 305 AND Y = 119 else
"110111011111" when X = 306 AND Y = 119 else
"110111011111" when X = 307 AND Y = 119 else
"110111011111" when X = 308 AND Y = 119 else
"110111011111" when X = 309 AND Y = 119 else
"110111011111" when X = 310 AND Y = 119 else
"110111011111" when X = 311 AND Y = 119 else
"110111011111" when X = 312 AND Y = 119 else
"110111011111" when X = 313 AND Y = 119 else
"110111011111" when X = 314 AND Y = 119 else
"110111011111" when X = 315 AND Y = 119 else
"110111011111" when X = 316 AND Y = 119 else
"110111011111" when X = 317 AND Y = 119 else
"110111011111" when X = 318 AND Y = 119 else
"110111011111" when X = 319 AND Y = 119 else
"110111011111" when X = 320 AND Y = 119 else
"110111011111" when X = 321 AND Y = 119 else
"110111011111" when X = 322 AND Y = 119 else
"110111011111" when X = 323 AND Y = 119 else
"110111011111" when X = 324 AND Y = 119 else
"100010011101" when X = 0 AND Y = 120 else
"100010011101" when X = 1 AND Y = 120 else
"100010011101" when X = 2 AND Y = 120 else
"100010011101" when X = 3 AND Y = 120 else
"100010011101" when X = 4 AND Y = 120 else
"100010011101" when X = 5 AND Y = 120 else
"100010011101" when X = 6 AND Y = 120 else
"100010011101" when X = 7 AND Y = 120 else
"100010011101" when X = 8 AND Y = 120 else
"100010011101" when X = 9 AND Y = 120 else
"100010011101" when X = 10 AND Y = 120 else
"100010011101" when X = 11 AND Y = 120 else
"100010011101" when X = 12 AND Y = 120 else
"100010011101" when X = 13 AND Y = 120 else
"100010011101" when X = 14 AND Y = 120 else
"100010011101" when X = 15 AND Y = 120 else
"100010011101" when X = 16 AND Y = 120 else
"100010011101" when X = 17 AND Y = 120 else
"100010011101" when X = 18 AND Y = 120 else
"100010011101" when X = 19 AND Y = 120 else
"100010011101" when X = 20 AND Y = 120 else
"100010011101" when X = 21 AND Y = 120 else
"100010011101" when X = 22 AND Y = 120 else
"100010011101" when X = 23 AND Y = 120 else
"100010011101" when X = 24 AND Y = 120 else
"100010011101" when X = 25 AND Y = 120 else
"100010011101" when X = 26 AND Y = 120 else
"100010011101" when X = 27 AND Y = 120 else
"100010011101" when X = 28 AND Y = 120 else
"100010011101" when X = 29 AND Y = 120 else
"100010011101" when X = 30 AND Y = 120 else
"100010011101" when X = 31 AND Y = 120 else
"100010011101" when X = 32 AND Y = 120 else
"100010011101" when X = 33 AND Y = 120 else
"100010011101" when X = 34 AND Y = 120 else
"100010011101" when X = 35 AND Y = 120 else
"100010011101" when X = 36 AND Y = 120 else
"100010011101" when X = 37 AND Y = 120 else
"100010011101" when X = 38 AND Y = 120 else
"100010011101" when X = 39 AND Y = 120 else
"110111011111" when X = 40 AND Y = 120 else
"110111011111" when X = 41 AND Y = 120 else
"110111011111" when X = 42 AND Y = 120 else
"110111011111" when X = 43 AND Y = 120 else
"110111011111" when X = 44 AND Y = 120 else
"110111011111" when X = 45 AND Y = 120 else
"110111011111" when X = 46 AND Y = 120 else
"110111011111" when X = 47 AND Y = 120 else
"110111011111" when X = 48 AND Y = 120 else
"110111011111" when X = 49 AND Y = 120 else
"110111011111" when X = 50 AND Y = 120 else
"110111011111" when X = 51 AND Y = 120 else
"110111011111" when X = 52 AND Y = 120 else
"110111011111" when X = 53 AND Y = 120 else
"110111011111" when X = 54 AND Y = 120 else
"110111011111" when X = 55 AND Y = 120 else
"110111011111" when X = 56 AND Y = 120 else
"110111011111" when X = 57 AND Y = 120 else
"110111011111" when X = 58 AND Y = 120 else
"110111011111" when X = 59 AND Y = 120 else
"110111011111" when X = 60 AND Y = 120 else
"110111011111" when X = 61 AND Y = 120 else
"110111011111" when X = 62 AND Y = 120 else
"110111011111" when X = 63 AND Y = 120 else
"110111011111" when X = 64 AND Y = 120 else
"110111011111" when X = 65 AND Y = 120 else
"110111011111" when X = 66 AND Y = 120 else
"110111011111" when X = 67 AND Y = 120 else
"110111011111" when X = 68 AND Y = 120 else
"110111011111" when X = 69 AND Y = 120 else
"110111011111" when X = 70 AND Y = 120 else
"110111011111" when X = 71 AND Y = 120 else
"110111011111" when X = 72 AND Y = 120 else
"110111011111" when X = 73 AND Y = 120 else
"110111011111" when X = 74 AND Y = 120 else
"110111011111" when X = 75 AND Y = 120 else
"110111011111" when X = 76 AND Y = 120 else
"110111011111" when X = 77 AND Y = 120 else
"110111011111" when X = 78 AND Y = 120 else
"110111011111" when X = 79 AND Y = 120 else
"110111011111" when X = 80 AND Y = 120 else
"110111011111" when X = 81 AND Y = 120 else
"110111011111" when X = 82 AND Y = 120 else
"110111011111" when X = 83 AND Y = 120 else
"110111011111" when X = 84 AND Y = 120 else
"110111011111" when X = 85 AND Y = 120 else
"110111011111" when X = 86 AND Y = 120 else
"110111011111" when X = 87 AND Y = 120 else
"110111011111" when X = 88 AND Y = 120 else
"110111011111" when X = 89 AND Y = 120 else
"110111011111" when X = 90 AND Y = 120 else
"110111011111" when X = 91 AND Y = 120 else
"110111011111" when X = 92 AND Y = 120 else
"110111011111" when X = 93 AND Y = 120 else
"110111011111" when X = 94 AND Y = 120 else
"110111011111" when X = 95 AND Y = 120 else
"110111011111" when X = 96 AND Y = 120 else
"110111011111" when X = 97 AND Y = 120 else
"110111011111" when X = 98 AND Y = 120 else
"110111011111" when X = 99 AND Y = 120 else
"110111011111" when X = 100 AND Y = 120 else
"110111011111" when X = 101 AND Y = 120 else
"110111011111" when X = 102 AND Y = 120 else
"110111011111" when X = 103 AND Y = 120 else
"110111011111" when X = 104 AND Y = 120 else
"110111011111" when X = 105 AND Y = 120 else
"110111011111" when X = 106 AND Y = 120 else
"110111011111" when X = 107 AND Y = 120 else
"110111011111" when X = 108 AND Y = 120 else
"110111011111" when X = 109 AND Y = 120 else
"110111011111" when X = 110 AND Y = 120 else
"110111011111" when X = 111 AND Y = 120 else
"110111011111" when X = 112 AND Y = 120 else
"110111011111" when X = 113 AND Y = 120 else
"110111011111" when X = 114 AND Y = 120 else
"110111011111" when X = 115 AND Y = 120 else
"110111011111" when X = 116 AND Y = 120 else
"110111011111" when X = 117 AND Y = 120 else
"110111011111" when X = 118 AND Y = 120 else
"110111011111" when X = 119 AND Y = 120 else
"110111011111" when X = 120 AND Y = 120 else
"110111011111" when X = 121 AND Y = 120 else
"110111011111" when X = 122 AND Y = 120 else
"110111011111" when X = 123 AND Y = 120 else
"110111011111" when X = 124 AND Y = 120 else
"110111011111" when X = 125 AND Y = 120 else
"110111011111" when X = 126 AND Y = 120 else
"110111011111" when X = 127 AND Y = 120 else
"110111011111" when X = 128 AND Y = 120 else
"110111011111" when X = 129 AND Y = 120 else
"110111011111" when X = 130 AND Y = 120 else
"110111011111" when X = 131 AND Y = 120 else
"110111011111" when X = 132 AND Y = 120 else
"110111011111" when X = 133 AND Y = 120 else
"110111011111" when X = 134 AND Y = 120 else
"110111011111" when X = 135 AND Y = 120 else
"110111011111" when X = 136 AND Y = 120 else
"110111011111" when X = 137 AND Y = 120 else
"110111011111" when X = 138 AND Y = 120 else
"110111011111" when X = 139 AND Y = 120 else
"110111011111" when X = 140 AND Y = 120 else
"110111011111" when X = 141 AND Y = 120 else
"110111011111" when X = 142 AND Y = 120 else
"110111011111" when X = 143 AND Y = 120 else
"110111011111" when X = 144 AND Y = 120 else
"110111011111" when X = 145 AND Y = 120 else
"110111011111" when X = 146 AND Y = 120 else
"110111011111" when X = 147 AND Y = 120 else
"110111011111" when X = 148 AND Y = 120 else
"110111011111" when X = 149 AND Y = 120 else
"110111011111" when X = 150 AND Y = 120 else
"110111011111" when X = 151 AND Y = 120 else
"110111011111" when X = 152 AND Y = 120 else
"110111011111" when X = 153 AND Y = 120 else
"110111011111" when X = 154 AND Y = 120 else
"110111011111" when X = 155 AND Y = 120 else
"110111011111" when X = 156 AND Y = 120 else
"110111011111" when X = 157 AND Y = 120 else
"110111011111" when X = 158 AND Y = 120 else
"110111011111" when X = 159 AND Y = 120 else
"110111011111" when X = 160 AND Y = 120 else
"110111011111" when X = 161 AND Y = 120 else
"110111011111" when X = 162 AND Y = 120 else
"110111011111" when X = 163 AND Y = 120 else
"110111011111" when X = 164 AND Y = 120 else
"111111111111" when X = 165 AND Y = 120 else
"111111111111" when X = 166 AND Y = 120 else
"111111111111" when X = 167 AND Y = 120 else
"111111111111" when X = 168 AND Y = 120 else
"111111111111" when X = 169 AND Y = 120 else
"111111111111" when X = 170 AND Y = 120 else
"111111111111" when X = 171 AND Y = 120 else
"111111111111" when X = 172 AND Y = 120 else
"111111111111" when X = 173 AND Y = 120 else
"111111111111" when X = 174 AND Y = 120 else
"111111111111" when X = 175 AND Y = 120 else
"111111111111" when X = 176 AND Y = 120 else
"111111111111" when X = 177 AND Y = 120 else
"111111111111" when X = 178 AND Y = 120 else
"111111111111" when X = 179 AND Y = 120 else
"111111111111" when X = 180 AND Y = 120 else
"111111111111" when X = 181 AND Y = 120 else
"111111111111" when X = 182 AND Y = 120 else
"111111111111" when X = 183 AND Y = 120 else
"111111111111" when X = 184 AND Y = 120 else
"111111111111" when X = 185 AND Y = 120 else
"111111111111" when X = 186 AND Y = 120 else
"111111111111" when X = 187 AND Y = 120 else
"111111111111" when X = 188 AND Y = 120 else
"111111111111" when X = 189 AND Y = 120 else
"110111011111" when X = 190 AND Y = 120 else
"110111011111" when X = 191 AND Y = 120 else
"110111011111" when X = 192 AND Y = 120 else
"110111011111" when X = 193 AND Y = 120 else
"110111011111" when X = 194 AND Y = 120 else
"110111011111" when X = 195 AND Y = 120 else
"110111011111" when X = 196 AND Y = 120 else
"110111011111" when X = 197 AND Y = 120 else
"110111011111" when X = 198 AND Y = 120 else
"110111011111" when X = 199 AND Y = 120 else
"110111011111" when X = 200 AND Y = 120 else
"110111011111" when X = 201 AND Y = 120 else
"110111011111" when X = 202 AND Y = 120 else
"110111011111" when X = 203 AND Y = 120 else
"110111011111" when X = 204 AND Y = 120 else
"110111011111" when X = 205 AND Y = 120 else
"110111011111" when X = 206 AND Y = 120 else
"110111011111" when X = 207 AND Y = 120 else
"110111011111" when X = 208 AND Y = 120 else
"110111011111" when X = 209 AND Y = 120 else
"110111011111" when X = 210 AND Y = 120 else
"110111011111" when X = 211 AND Y = 120 else
"110111011111" when X = 212 AND Y = 120 else
"110111011111" when X = 213 AND Y = 120 else
"110111011111" when X = 214 AND Y = 120 else
"110111011111" when X = 215 AND Y = 120 else
"110111011111" when X = 216 AND Y = 120 else
"110111011111" when X = 217 AND Y = 120 else
"110111011111" when X = 218 AND Y = 120 else
"110111011111" when X = 219 AND Y = 120 else
"110111011111" when X = 220 AND Y = 120 else
"110111011111" when X = 221 AND Y = 120 else
"110111011111" when X = 222 AND Y = 120 else
"110111011111" when X = 223 AND Y = 120 else
"110111011111" when X = 224 AND Y = 120 else
"110111011111" when X = 225 AND Y = 120 else
"110111011111" when X = 226 AND Y = 120 else
"110111011111" when X = 227 AND Y = 120 else
"110111011111" when X = 228 AND Y = 120 else
"110111011111" when X = 229 AND Y = 120 else
"110111011111" when X = 230 AND Y = 120 else
"110111011111" when X = 231 AND Y = 120 else
"110111011111" when X = 232 AND Y = 120 else
"110111011111" when X = 233 AND Y = 120 else
"110111011111" when X = 234 AND Y = 120 else
"110111011111" when X = 235 AND Y = 120 else
"110111011111" when X = 236 AND Y = 120 else
"110111011111" when X = 237 AND Y = 120 else
"110111011111" when X = 238 AND Y = 120 else
"110111011111" when X = 239 AND Y = 120 else
"110111011111" when X = 240 AND Y = 120 else
"110111011111" when X = 241 AND Y = 120 else
"110111011111" when X = 242 AND Y = 120 else
"110111011111" when X = 243 AND Y = 120 else
"110111011111" when X = 244 AND Y = 120 else
"110111011111" when X = 245 AND Y = 120 else
"110111011111" when X = 246 AND Y = 120 else
"110111011111" when X = 247 AND Y = 120 else
"110111011111" when X = 248 AND Y = 120 else
"110111011111" when X = 249 AND Y = 120 else
"110111011111" when X = 250 AND Y = 120 else
"110111011111" when X = 251 AND Y = 120 else
"110111011111" when X = 252 AND Y = 120 else
"110111011111" when X = 253 AND Y = 120 else
"110111011111" when X = 254 AND Y = 120 else
"110111011111" when X = 255 AND Y = 120 else
"110111011111" when X = 256 AND Y = 120 else
"110111011111" when X = 257 AND Y = 120 else
"110111011111" when X = 258 AND Y = 120 else
"110111011111" when X = 259 AND Y = 120 else
"110111011111" when X = 260 AND Y = 120 else
"110111011111" when X = 261 AND Y = 120 else
"110111011111" when X = 262 AND Y = 120 else
"110111011111" when X = 263 AND Y = 120 else
"110111011111" when X = 264 AND Y = 120 else
"110111011111" when X = 265 AND Y = 120 else
"110111011111" when X = 266 AND Y = 120 else
"110111011111" when X = 267 AND Y = 120 else
"110111011111" when X = 268 AND Y = 120 else
"110111011111" when X = 269 AND Y = 120 else
"110111011111" when X = 270 AND Y = 120 else
"110111011111" when X = 271 AND Y = 120 else
"110111011111" when X = 272 AND Y = 120 else
"110111011111" when X = 273 AND Y = 120 else
"110111011111" when X = 274 AND Y = 120 else
"110111011111" when X = 275 AND Y = 120 else
"110111011111" when X = 276 AND Y = 120 else
"110111011111" when X = 277 AND Y = 120 else
"110111011111" when X = 278 AND Y = 120 else
"110111011111" when X = 279 AND Y = 120 else
"110111011111" when X = 280 AND Y = 120 else
"110111011111" when X = 281 AND Y = 120 else
"110111011111" when X = 282 AND Y = 120 else
"110111011111" when X = 283 AND Y = 120 else
"110111011111" when X = 284 AND Y = 120 else
"110111011111" when X = 285 AND Y = 120 else
"110111011111" when X = 286 AND Y = 120 else
"110111011111" when X = 287 AND Y = 120 else
"110111011111" when X = 288 AND Y = 120 else
"110111011111" when X = 289 AND Y = 120 else
"110111011111" when X = 290 AND Y = 120 else
"110111011111" when X = 291 AND Y = 120 else
"110111011111" when X = 292 AND Y = 120 else
"110111011111" when X = 293 AND Y = 120 else
"110111011111" when X = 294 AND Y = 120 else
"110111011111" when X = 295 AND Y = 120 else
"110111011111" when X = 296 AND Y = 120 else
"110111011111" when X = 297 AND Y = 120 else
"110111011111" when X = 298 AND Y = 120 else
"110111011111" when X = 299 AND Y = 120 else
"110111011111" when X = 300 AND Y = 120 else
"110111011111" when X = 301 AND Y = 120 else
"110111011111" when X = 302 AND Y = 120 else
"110111011111" when X = 303 AND Y = 120 else
"110111011111" when X = 304 AND Y = 120 else
"110111011111" when X = 305 AND Y = 120 else
"110111011111" when X = 306 AND Y = 120 else
"110111011111" when X = 307 AND Y = 120 else
"110111011111" when X = 308 AND Y = 120 else
"110111011111" when X = 309 AND Y = 120 else
"110111011111" when X = 310 AND Y = 120 else
"110111011111" when X = 311 AND Y = 120 else
"110111011111" when X = 312 AND Y = 120 else
"110111011111" when X = 313 AND Y = 120 else
"110111011111" when X = 314 AND Y = 120 else
"110111011111" when X = 315 AND Y = 120 else
"110111011111" when X = 316 AND Y = 120 else
"110111011111" when X = 317 AND Y = 120 else
"110111011111" when X = 318 AND Y = 120 else
"110111011111" when X = 319 AND Y = 120 else
"110111011111" when X = 320 AND Y = 120 else
"110111011111" when X = 321 AND Y = 120 else
"110111011111" when X = 322 AND Y = 120 else
"110111011111" when X = 323 AND Y = 120 else
"110111011111" when X = 324 AND Y = 120 else
"100010011101" when X = 0 AND Y = 121 else
"100010011101" when X = 1 AND Y = 121 else
"100010011101" when X = 2 AND Y = 121 else
"100010011101" when X = 3 AND Y = 121 else
"100010011101" when X = 4 AND Y = 121 else
"100010011101" when X = 5 AND Y = 121 else
"100010011101" when X = 6 AND Y = 121 else
"100010011101" when X = 7 AND Y = 121 else
"100010011101" when X = 8 AND Y = 121 else
"100010011101" when X = 9 AND Y = 121 else
"100010011101" when X = 10 AND Y = 121 else
"100010011101" when X = 11 AND Y = 121 else
"100010011101" when X = 12 AND Y = 121 else
"100010011101" when X = 13 AND Y = 121 else
"100010011101" when X = 14 AND Y = 121 else
"100010011101" when X = 15 AND Y = 121 else
"100010011101" when X = 16 AND Y = 121 else
"100010011101" when X = 17 AND Y = 121 else
"100010011101" when X = 18 AND Y = 121 else
"100010011101" when X = 19 AND Y = 121 else
"100010011101" when X = 20 AND Y = 121 else
"100010011101" when X = 21 AND Y = 121 else
"100010011101" when X = 22 AND Y = 121 else
"100010011101" when X = 23 AND Y = 121 else
"100010011101" when X = 24 AND Y = 121 else
"100010011101" when X = 25 AND Y = 121 else
"100010011101" when X = 26 AND Y = 121 else
"100010011101" when X = 27 AND Y = 121 else
"100010011101" when X = 28 AND Y = 121 else
"100010011101" when X = 29 AND Y = 121 else
"100010011101" when X = 30 AND Y = 121 else
"100010011101" when X = 31 AND Y = 121 else
"100010011101" when X = 32 AND Y = 121 else
"100010011101" when X = 33 AND Y = 121 else
"100010011101" when X = 34 AND Y = 121 else
"100010011101" when X = 35 AND Y = 121 else
"100010011101" when X = 36 AND Y = 121 else
"100010011101" when X = 37 AND Y = 121 else
"100010011101" when X = 38 AND Y = 121 else
"100010011101" when X = 39 AND Y = 121 else
"110111011111" when X = 40 AND Y = 121 else
"110111011111" when X = 41 AND Y = 121 else
"110111011111" when X = 42 AND Y = 121 else
"110111011111" when X = 43 AND Y = 121 else
"110111011111" when X = 44 AND Y = 121 else
"110111011111" when X = 45 AND Y = 121 else
"110111011111" when X = 46 AND Y = 121 else
"110111011111" when X = 47 AND Y = 121 else
"110111011111" when X = 48 AND Y = 121 else
"110111011111" when X = 49 AND Y = 121 else
"110111011111" when X = 50 AND Y = 121 else
"110111011111" when X = 51 AND Y = 121 else
"110111011111" when X = 52 AND Y = 121 else
"110111011111" when X = 53 AND Y = 121 else
"110111011111" when X = 54 AND Y = 121 else
"110111011111" when X = 55 AND Y = 121 else
"110111011111" when X = 56 AND Y = 121 else
"110111011111" when X = 57 AND Y = 121 else
"110111011111" when X = 58 AND Y = 121 else
"110111011111" when X = 59 AND Y = 121 else
"110111011111" when X = 60 AND Y = 121 else
"110111011111" when X = 61 AND Y = 121 else
"110111011111" when X = 62 AND Y = 121 else
"110111011111" when X = 63 AND Y = 121 else
"110111011111" when X = 64 AND Y = 121 else
"110111011111" when X = 65 AND Y = 121 else
"110111011111" when X = 66 AND Y = 121 else
"110111011111" when X = 67 AND Y = 121 else
"110111011111" when X = 68 AND Y = 121 else
"110111011111" when X = 69 AND Y = 121 else
"110111011111" when X = 70 AND Y = 121 else
"110111011111" when X = 71 AND Y = 121 else
"110111011111" when X = 72 AND Y = 121 else
"110111011111" when X = 73 AND Y = 121 else
"110111011111" when X = 74 AND Y = 121 else
"110111011111" when X = 75 AND Y = 121 else
"110111011111" when X = 76 AND Y = 121 else
"110111011111" when X = 77 AND Y = 121 else
"110111011111" when X = 78 AND Y = 121 else
"110111011111" when X = 79 AND Y = 121 else
"110111011111" when X = 80 AND Y = 121 else
"110111011111" when X = 81 AND Y = 121 else
"110111011111" when X = 82 AND Y = 121 else
"110111011111" when X = 83 AND Y = 121 else
"110111011111" when X = 84 AND Y = 121 else
"110111011111" when X = 85 AND Y = 121 else
"110111011111" when X = 86 AND Y = 121 else
"110111011111" when X = 87 AND Y = 121 else
"110111011111" when X = 88 AND Y = 121 else
"110111011111" when X = 89 AND Y = 121 else
"110111011111" when X = 90 AND Y = 121 else
"110111011111" when X = 91 AND Y = 121 else
"110111011111" when X = 92 AND Y = 121 else
"110111011111" when X = 93 AND Y = 121 else
"110111011111" when X = 94 AND Y = 121 else
"110111011111" when X = 95 AND Y = 121 else
"110111011111" when X = 96 AND Y = 121 else
"110111011111" when X = 97 AND Y = 121 else
"110111011111" when X = 98 AND Y = 121 else
"110111011111" when X = 99 AND Y = 121 else
"110111011111" when X = 100 AND Y = 121 else
"110111011111" when X = 101 AND Y = 121 else
"110111011111" when X = 102 AND Y = 121 else
"110111011111" when X = 103 AND Y = 121 else
"110111011111" when X = 104 AND Y = 121 else
"110111011111" when X = 105 AND Y = 121 else
"110111011111" when X = 106 AND Y = 121 else
"110111011111" when X = 107 AND Y = 121 else
"110111011111" when X = 108 AND Y = 121 else
"110111011111" when X = 109 AND Y = 121 else
"110111011111" when X = 110 AND Y = 121 else
"110111011111" when X = 111 AND Y = 121 else
"110111011111" when X = 112 AND Y = 121 else
"110111011111" when X = 113 AND Y = 121 else
"110111011111" when X = 114 AND Y = 121 else
"110111011111" when X = 115 AND Y = 121 else
"110111011111" when X = 116 AND Y = 121 else
"110111011111" when X = 117 AND Y = 121 else
"110111011111" when X = 118 AND Y = 121 else
"110111011111" when X = 119 AND Y = 121 else
"110111011111" when X = 120 AND Y = 121 else
"110111011111" when X = 121 AND Y = 121 else
"110111011111" when X = 122 AND Y = 121 else
"110111011111" when X = 123 AND Y = 121 else
"110111011111" when X = 124 AND Y = 121 else
"110111011111" when X = 125 AND Y = 121 else
"110111011111" when X = 126 AND Y = 121 else
"110111011111" when X = 127 AND Y = 121 else
"110111011111" when X = 128 AND Y = 121 else
"110111011111" when X = 129 AND Y = 121 else
"110111011111" when X = 130 AND Y = 121 else
"110111011111" when X = 131 AND Y = 121 else
"110111011111" when X = 132 AND Y = 121 else
"110111011111" when X = 133 AND Y = 121 else
"110111011111" when X = 134 AND Y = 121 else
"110111011111" when X = 135 AND Y = 121 else
"110111011111" when X = 136 AND Y = 121 else
"110111011111" when X = 137 AND Y = 121 else
"110111011111" when X = 138 AND Y = 121 else
"110111011111" when X = 139 AND Y = 121 else
"110111011111" when X = 140 AND Y = 121 else
"110111011111" when X = 141 AND Y = 121 else
"110111011111" when X = 142 AND Y = 121 else
"110111011111" when X = 143 AND Y = 121 else
"110111011111" when X = 144 AND Y = 121 else
"110111011111" when X = 145 AND Y = 121 else
"110111011111" when X = 146 AND Y = 121 else
"110111011111" when X = 147 AND Y = 121 else
"110111011111" when X = 148 AND Y = 121 else
"110111011111" when X = 149 AND Y = 121 else
"110111011111" when X = 150 AND Y = 121 else
"110111011111" when X = 151 AND Y = 121 else
"110111011111" when X = 152 AND Y = 121 else
"110111011111" when X = 153 AND Y = 121 else
"110111011111" when X = 154 AND Y = 121 else
"110111011111" when X = 155 AND Y = 121 else
"110111011111" when X = 156 AND Y = 121 else
"110111011111" when X = 157 AND Y = 121 else
"110111011111" when X = 158 AND Y = 121 else
"110111011111" when X = 159 AND Y = 121 else
"110111011111" when X = 160 AND Y = 121 else
"110111011111" when X = 161 AND Y = 121 else
"110111011111" when X = 162 AND Y = 121 else
"110111011111" when X = 163 AND Y = 121 else
"110111011111" when X = 164 AND Y = 121 else
"111111111111" when X = 165 AND Y = 121 else
"111111111111" when X = 166 AND Y = 121 else
"111111111111" when X = 167 AND Y = 121 else
"111111111111" when X = 168 AND Y = 121 else
"111111111111" when X = 169 AND Y = 121 else
"111111111111" when X = 170 AND Y = 121 else
"111111111111" when X = 171 AND Y = 121 else
"111111111111" when X = 172 AND Y = 121 else
"111111111111" when X = 173 AND Y = 121 else
"111111111111" when X = 174 AND Y = 121 else
"111111111111" when X = 175 AND Y = 121 else
"111111111111" when X = 176 AND Y = 121 else
"111111111111" when X = 177 AND Y = 121 else
"111111111111" when X = 178 AND Y = 121 else
"111111111111" when X = 179 AND Y = 121 else
"111111111111" when X = 180 AND Y = 121 else
"111111111111" when X = 181 AND Y = 121 else
"111111111111" when X = 182 AND Y = 121 else
"111111111111" when X = 183 AND Y = 121 else
"111111111111" when X = 184 AND Y = 121 else
"111111111111" when X = 185 AND Y = 121 else
"111111111111" when X = 186 AND Y = 121 else
"111111111111" when X = 187 AND Y = 121 else
"111111111111" when X = 188 AND Y = 121 else
"111111111111" when X = 189 AND Y = 121 else
"110111011111" when X = 190 AND Y = 121 else
"110111011111" when X = 191 AND Y = 121 else
"110111011111" when X = 192 AND Y = 121 else
"110111011111" when X = 193 AND Y = 121 else
"110111011111" when X = 194 AND Y = 121 else
"110111011111" when X = 195 AND Y = 121 else
"110111011111" when X = 196 AND Y = 121 else
"110111011111" when X = 197 AND Y = 121 else
"110111011111" when X = 198 AND Y = 121 else
"110111011111" when X = 199 AND Y = 121 else
"110111011111" when X = 200 AND Y = 121 else
"110111011111" when X = 201 AND Y = 121 else
"110111011111" when X = 202 AND Y = 121 else
"110111011111" when X = 203 AND Y = 121 else
"110111011111" when X = 204 AND Y = 121 else
"110111011111" when X = 205 AND Y = 121 else
"110111011111" when X = 206 AND Y = 121 else
"110111011111" when X = 207 AND Y = 121 else
"110111011111" when X = 208 AND Y = 121 else
"110111011111" when X = 209 AND Y = 121 else
"110111011111" when X = 210 AND Y = 121 else
"110111011111" when X = 211 AND Y = 121 else
"110111011111" when X = 212 AND Y = 121 else
"110111011111" when X = 213 AND Y = 121 else
"110111011111" when X = 214 AND Y = 121 else
"110111011111" when X = 215 AND Y = 121 else
"110111011111" when X = 216 AND Y = 121 else
"110111011111" when X = 217 AND Y = 121 else
"110111011111" when X = 218 AND Y = 121 else
"110111011111" when X = 219 AND Y = 121 else
"110111011111" when X = 220 AND Y = 121 else
"110111011111" when X = 221 AND Y = 121 else
"110111011111" when X = 222 AND Y = 121 else
"110111011111" when X = 223 AND Y = 121 else
"110111011111" when X = 224 AND Y = 121 else
"110111011111" when X = 225 AND Y = 121 else
"110111011111" when X = 226 AND Y = 121 else
"110111011111" when X = 227 AND Y = 121 else
"110111011111" when X = 228 AND Y = 121 else
"110111011111" when X = 229 AND Y = 121 else
"110111011111" when X = 230 AND Y = 121 else
"110111011111" when X = 231 AND Y = 121 else
"110111011111" when X = 232 AND Y = 121 else
"110111011111" when X = 233 AND Y = 121 else
"110111011111" when X = 234 AND Y = 121 else
"110111011111" when X = 235 AND Y = 121 else
"110111011111" when X = 236 AND Y = 121 else
"110111011111" when X = 237 AND Y = 121 else
"110111011111" when X = 238 AND Y = 121 else
"110111011111" when X = 239 AND Y = 121 else
"110111011111" when X = 240 AND Y = 121 else
"110111011111" when X = 241 AND Y = 121 else
"110111011111" when X = 242 AND Y = 121 else
"110111011111" when X = 243 AND Y = 121 else
"110111011111" when X = 244 AND Y = 121 else
"110111011111" when X = 245 AND Y = 121 else
"110111011111" when X = 246 AND Y = 121 else
"110111011111" when X = 247 AND Y = 121 else
"110111011111" when X = 248 AND Y = 121 else
"110111011111" when X = 249 AND Y = 121 else
"110111011111" when X = 250 AND Y = 121 else
"110111011111" when X = 251 AND Y = 121 else
"110111011111" when X = 252 AND Y = 121 else
"110111011111" when X = 253 AND Y = 121 else
"110111011111" when X = 254 AND Y = 121 else
"110111011111" when X = 255 AND Y = 121 else
"110111011111" when X = 256 AND Y = 121 else
"110111011111" when X = 257 AND Y = 121 else
"110111011111" when X = 258 AND Y = 121 else
"110111011111" when X = 259 AND Y = 121 else
"110111011111" when X = 260 AND Y = 121 else
"110111011111" when X = 261 AND Y = 121 else
"110111011111" when X = 262 AND Y = 121 else
"110111011111" when X = 263 AND Y = 121 else
"110111011111" when X = 264 AND Y = 121 else
"110111011111" when X = 265 AND Y = 121 else
"110111011111" when X = 266 AND Y = 121 else
"110111011111" when X = 267 AND Y = 121 else
"110111011111" when X = 268 AND Y = 121 else
"110111011111" when X = 269 AND Y = 121 else
"110111011111" when X = 270 AND Y = 121 else
"110111011111" when X = 271 AND Y = 121 else
"110111011111" when X = 272 AND Y = 121 else
"110111011111" when X = 273 AND Y = 121 else
"110111011111" when X = 274 AND Y = 121 else
"110111011111" when X = 275 AND Y = 121 else
"110111011111" when X = 276 AND Y = 121 else
"110111011111" when X = 277 AND Y = 121 else
"110111011111" when X = 278 AND Y = 121 else
"110111011111" when X = 279 AND Y = 121 else
"110111011111" when X = 280 AND Y = 121 else
"110111011111" when X = 281 AND Y = 121 else
"110111011111" when X = 282 AND Y = 121 else
"110111011111" when X = 283 AND Y = 121 else
"110111011111" when X = 284 AND Y = 121 else
"110111011111" when X = 285 AND Y = 121 else
"110111011111" when X = 286 AND Y = 121 else
"110111011111" when X = 287 AND Y = 121 else
"110111011111" when X = 288 AND Y = 121 else
"110111011111" when X = 289 AND Y = 121 else
"110111011111" when X = 290 AND Y = 121 else
"110111011111" when X = 291 AND Y = 121 else
"110111011111" when X = 292 AND Y = 121 else
"110111011111" when X = 293 AND Y = 121 else
"110111011111" when X = 294 AND Y = 121 else
"110111011111" when X = 295 AND Y = 121 else
"110111011111" when X = 296 AND Y = 121 else
"110111011111" when X = 297 AND Y = 121 else
"110111011111" when X = 298 AND Y = 121 else
"110111011111" when X = 299 AND Y = 121 else
"110111011111" when X = 300 AND Y = 121 else
"110111011111" when X = 301 AND Y = 121 else
"110111011111" when X = 302 AND Y = 121 else
"110111011111" when X = 303 AND Y = 121 else
"110111011111" when X = 304 AND Y = 121 else
"110111011111" when X = 305 AND Y = 121 else
"110111011111" when X = 306 AND Y = 121 else
"110111011111" when X = 307 AND Y = 121 else
"110111011111" when X = 308 AND Y = 121 else
"110111011111" when X = 309 AND Y = 121 else
"110111011111" when X = 310 AND Y = 121 else
"110111011111" when X = 311 AND Y = 121 else
"110111011111" when X = 312 AND Y = 121 else
"110111011111" when X = 313 AND Y = 121 else
"110111011111" when X = 314 AND Y = 121 else
"110111011111" when X = 315 AND Y = 121 else
"110111011111" when X = 316 AND Y = 121 else
"110111011111" when X = 317 AND Y = 121 else
"110111011111" when X = 318 AND Y = 121 else
"110111011111" when X = 319 AND Y = 121 else
"110111011111" when X = 320 AND Y = 121 else
"110111011111" when X = 321 AND Y = 121 else
"110111011111" when X = 322 AND Y = 121 else
"110111011111" when X = 323 AND Y = 121 else
"110111011111" when X = 324 AND Y = 121 else
"100010011101" when X = 0 AND Y = 122 else
"100010011101" when X = 1 AND Y = 122 else
"100010011101" when X = 2 AND Y = 122 else
"100010011101" when X = 3 AND Y = 122 else
"100010011101" when X = 4 AND Y = 122 else
"100010011101" when X = 5 AND Y = 122 else
"100010011101" when X = 6 AND Y = 122 else
"100010011101" when X = 7 AND Y = 122 else
"100010011101" when X = 8 AND Y = 122 else
"100010011101" when X = 9 AND Y = 122 else
"100010011101" when X = 10 AND Y = 122 else
"100010011101" when X = 11 AND Y = 122 else
"100010011101" when X = 12 AND Y = 122 else
"100010011101" when X = 13 AND Y = 122 else
"100010011101" when X = 14 AND Y = 122 else
"100010011101" when X = 15 AND Y = 122 else
"100010011101" when X = 16 AND Y = 122 else
"100010011101" when X = 17 AND Y = 122 else
"100010011101" when X = 18 AND Y = 122 else
"100010011101" when X = 19 AND Y = 122 else
"100010011101" when X = 20 AND Y = 122 else
"100010011101" when X = 21 AND Y = 122 else
"100010011101" when X = 22 AND Y = 122 else
"100010011101" when X = 23 AND Y = 122 else
"100010011101" when X = 24 AND Y = 122 else
"100010011101" when X = 25 AND Y = 122 else
"100010011101" when X = 26 AND Y = 122 else
"100010011101" when X = 27 AND Y = 122 else
"100010011101" when X = 28 AND Y = 122 else
"100010011101" when X = 29 AND Y = 122 else
"100010011101" when X = 30 AND Y = 122 else
"100010011101" when X = 31 AND Y = 122 else
"100010011101" when X = 32 AND Y = 122 else
"100010011101" when X = 33 AND Y = 122 else
"100010011101" when X = 34 AND Y = 122 else
"100010011101" when X = 35 AND Y = 122 else
"100010011101" when X = 36 AND Y = 122 else
"100010011101" when X = 37 AND Y = 122 else
"100010011101" when X = 38 AND Y = 122 else
"100010011101" when X = 39 AND Y = 122 else
"110111011111" when X = 40 AND Y = 122 else
"110111011111" when X = 41 AND Y = 122 else
"110111011111" when X = 42 AND Y = 122 else
"110111011111" when X = 43 AND Y = 122 else
"110111011111" when X = 44 AND Y = 122 else
"110111011111" when X = 45 AND Y = 122 else
"110111011111" when X = 46 AND Y = 122 else
"110111011111" when X = 47 AND Y = 122 else
"110111011111" when X = 48 AND Y = 122 else
"110111011111" when X = 49 AND Y = 122 else
"110111011111" when X = 50 AND Y = 122 else
"110111011111" when X = 51 AND Y = 122 else
"110111011111" when X = 52 AND Y = 122 else
"110111011111" when X = 53 AND Y = 122 else
"110111011111" when X = 54 AND Y = 122 else
"110111011111" when X = 55 AND Y = 122 else
"110111011111" when X = 56 AND Y = 122 else
"110111011111" when X = 57 AND Y = 122 else
"110111011111" when X = 58 AND Y = 122 else
"110111011111" when X = 59 AND Y = 122 else
"110111011111" when X = 60 AND Y = 122 else
"110111011111" when X = 61 AND Y = 122 else
"110111011111" when X = 62 AND Y = 122 else
"110111011111" when X = 63 AND Y = 122 else
"110111011111" when X = 64 AND Y = 122 else
"110111011111" when X = 65 AND Y = 122 else
"110111011111" when X = 66 AND Y = 122 else
"110111011111" when X = 67 AND Y = 122 else
"110111011111" when X = 68 AND Y = 122 else
"110111011111" when X = 69 AND Y = 122 else
"110111011111" when X = 70 AND Y = 122 else
"110111011111" when X = 71 AND Y = 122 else
"110111011111" when X = 72 AND Y = 122 else
"110111011111" when X = 73 AND Y = 122 else
"110111011111" when X = 74 AND Y = 122 else
"110111011111" when X = 75 AND Y = 122 else
"110111011111" when X = 76 AND Y = 122 else
"110111011111" when X = 77 AND Y = 122 else
"110111011111" when X = 78 AND Y = 122 else
"110111011111" when X = 79 AND Y = 122 else
"110111011111" when X = 80 AND Y = 122 else
"110111011111" when X = 81 AND Y = 122 else
"110111011111" when X = 82 AND Y = 122 else
"110111011111" when X = 83 AND Y = 122 else
"110111011111" when X = 84 AND Y = 122 else
"110111011111" when X = 85 AND Y = 122 else
"110111011111" when X = 86 AND Y = 122 else
"110111011111" when X = 87 AND Y = 122 else
"110111011111" when X = 88 AND Y = 122 else
"110111011111" when X = 89 AND Y = 122 else
"110111011111" when X = 90 AND Y = 122 else
"110111011111" when X = 91 AND Y = 122 else
"110111011111" when X = 92 AND Y = 122 else
"110111011111" when X = 93 AND Y = 122 else
"110111011111" when X = 94 AND Y = 122 else
"110111011111" when X = 95 AND Y = 122 else
"110111011111" when X = 96 AND Y = 122 else
"110111011111" when X = 97 AND Y = 122 else
"110111011111" when X = 98 AND Y = 122 else
"110111011111" when X = 99 AND Y = 122 else
"110111011111" when X = 100 AND Y = 122 else
"110111011111" when X = 101 AND Y = 122 else
"110111011111" when X = 102 AND Y = 122 else
"110111011111" when X = 103 AND Y = 122 else
"110111011111" when X = 104 AND Y = 122 else
"110111011111" when X = 105 AND Y = 122 else
"110111011111" when X = 106 AND Y = 122 else
"110111011111" when X = 107 AND Y = 122 else
"110111011111" when X = 108 AND Y = 122 else
"110111011111" when X = 109 AND Y = 122 else
"110111011111" when X = 110 AND Y = 122 else
"110111011111" when X = 111 AND Y = 122 else
"110111011111" when X = 112 AND Y = 122 else
"110111011111" when X = 113 AND Y = 122 else
"110111011111" when X = 114 AND Y = 122 else
"110111011111" when X = 115 AND Y = 122 else
"110111011111" when X = 116 AND Y = 122 else
"110111011111" when X = 117 AND Y = 122 else
"110111011111" when X = 118 AND Y = 122 else
"110111011111" when X = 119 AND Y = 122 else
"110111011111" when X = 120 AND Y = 122 else
"110111011111" when X = 121 AND Y = 122 else
"110111011111" when X = 122 AND Y = 122 else
"110111011111" when X = 123 AND Y = 122 else
"110111011111" when X = 124 AND Y = 122 else
"110111011111" when X = 125 AND Y = 122 else
"110111011111" when X = 126 AND Y = 122 else
"110111011111" when X = 127 AND Y = 122 else
"110111011111" when X = 128 AND Y = 122 else
"110111011111" when X = 129 AND Y = 122 else
"110111011111" when X = 130 AND Y = 122 else
"110111011111" when X = 131 AND Y = 122 else
"110111011111" when X = 132 AND Y = 122 else
"110111011111" when X = 133 AND Y = 122 else
"110111011111" when X = 134 AND Y = 122 else
"110111011111" when X = 135 AND Y = 122 else
"110111011111" when X = 136 AND Y = 122 else
"110111011111" when X = 137 AND Y = 122 else
"110111011111" when X = 138 AND Y = 122 else
"110111011111" when X = 139 AND Y = 122 else
"110111011111" when X = 140 AND Y = 122 else
"110111011111" when X = 141 AND Y = 122 else
"110111011111" when X = 142 AND Y = 122 else
"110111011111" when X = 143 AND Y = 122 else
"110111011111" when X = 144 AND Y = 122 else
"110111011111" when X = 145 AND Y = 122 else
"110111011111" when X = 146 AND Y = 122 else
"110111011111" when X = 147 AND Y = 122 else
"110111011111" when X = 148 AND Y = 122 else
"110111011111" when X = 149 AND Y = 122 else
"110111011111" when X = 150 AND Y = 122 else
"110111011111" when X = 151 AND Y = 122 else
"110111011111" when X = 152 AND Y = 122 else
"110111011111" when X = 153 AND Y = 122 else
"110111011111" when X = 154 AND Y = 122 else
"110111011111" when X = 155 AND Y = 122 else
"110111011111" when X = 156 AND Y = 122 else
"110111011111" when X = 157 AND Y = 122 else
"110111011111" when X = 158 AND Y = 122 else
"110111011111" when X = 159 AND Y = 122 else
"110111011111" when X = 160 AND Y = 122 else
"110111011111" when X = 161 AND Y = 122 else
"110111011111" when X = 162 AND Y = 122 else
"110111011111" when X = 163 AND Y = 122 else
"110111011111" when X = 164 AND Y = 122 else
"111111111111" when X = 165 AND Y = 122 else
"111111111111" when X = 166 AND Y = 122 else
"111111111111" when X = 167 AND Y = 122 else
"111111111111" when X = 168 AND Y = 122 else
"111111111111" when X = 169 AND Y = 122 else
"111111111111" when X = 170 AND Y = 122 else
"111111111111" when X = 171 AND Y = 122 else
"111111111111" when X = 172 AND Y = 122 else
"111111111111" when X = 173 AND Y = 122 else
"111111111111" when X = 174 AND Y = 122 else
"111111111111" when X = 175 AND Y = 122 else
"111111111111" when X = 176 AND Y = 122 else
"111111111111" when X = 177 AND Y = 122 else
"111111111111" when X = 178 AND Y = 122 else
"111111111111" when X = 179 AND Y = 122 else
"111111111111" when X = 180 AND Y = 122 else
"111111111111" when X = 181 AND Y = 122 else
"111111111111" when X = 182 AND Y = 122 else
"111111111111" when X = 183 AND Y = 122 else
"111111111111" when X = 184 AND Y = 122 else
"111111111111" when X = 185 AND Y = 122 else
"111111111111" when X = 186 AND Y = 122 else
"111111111111" when X = 187 AND Y = 122 else
"111111111111" when X = 188 AND Y = 122 else
"111111111111" when X = 189 AND Y = 122 else
"110111011111" when X = 190 AND Y = 122 else
"110111011111" when X = 191 AND Y = 122 else
"110111011111" when X = 192 AND Y = 122 else
"110111011111" when X = 193 AND Y = 122 else
"110111011111" when X = 194 AND Y = 122 else
"110111011111" when X = 195 AND Y = 122 else
"110111011111" when X = 196 AND Y = 122 else
"110111011111" when X = 197 AND Y = 122 else
"110111011111" when X = 198 AND Y = 122 else
"110111011111" when X = 199 AND Y = 122 else
"110111011111" when X = 200 AND Y = 122 else
"110111011111" when X = 201 AND Y = 122 else
"110111011111" when X = 202 AND Y = 122 else
"110111011111" when X = 203 AND Y = 122 else
"110111011111" when X = 204 AND Y = 122 else
"110111011111" when X = 205 AND Y = 122 else
"110111011111" when X = 206 AND Y = 122 else
"110111011111" when X = 207 AND Y = 122 else
"110111011111" when X = 208 AND Y = 122 else
"110111011111" when X = 209 AND Y = 122 else
"110111011111" when X = 210 AND Y = 122 else
"110111011111" when X = 211 AND Y = 122 else
"110111011111" when X = 212 AND Y = 122 else
"110111011111" when X = 213 AND Y = 122 else
"110111011111" when X = 214 AND Y = 122 else
"110111011111" when X = 215 AND Y = 122 else
"110111011111" when X = 216 AND Y = 122 else
"110111011111" when X = 217 AND Y = 122 else
"110111011111" when X = 218 AND Y = 122 else
"110111011111" when X = 219 AND Y = 122 else
"110111011111" when X = 220 AND Y = 122 else
"110111011111" when X = 221 AND Y = 122 else
"110111011111" when X = 222 AND Y = 122 else
"110111011111" when X = 223 AND Y = 122 else
"110111011111" when X = 224 AND Y = 122 else
"110111011111" when X = 225 AND Y = 122 else
"110111011111" when X = 226 AND Y = 122 else
"110111011111" when X = 227 AND Y = 122 else
"110111011111" when X = 228 AND Y = 122 else
"110111011111" when X = 229 AND Y = 122 else
"110111011111" when X = 230 AND Y = 122 else
"110111011111" when X = 231 AND Y = 122 else
"110111011111" when X = 232 AND Y = 122 else
"110111011111" when X = 233 AND Y = 122 else
"110111011111" when X = 234 AND Y = 122 else
"110111011111" when X = 235 AND Y = 122 else
"110111011111" when X = 236 AND Y = 122 else
"110111011111" when X = 237 AND Y = 122 else
"110111011111" when X = 238 AND Y = 122 else
"110111011111" when X = 239 AND Y = 122 else
"110111011111" when X = 240 AND Y = 122 else
"110111011111" when X = 241 AND Y = 122 else
"110111011111" when X = 242 AND Y = 122 else
"110111011111" when X = 243 AND Y = 122 else
"110111011111" when X = 244 AND Y = 122 else
"110111011111" when X = 245 AND Y = 122 else
"110111011111" when X = 246 AND Y = 122 else
"110111011111" when X = 247 AND Y = 122 else
"110111011111" when X = 248 AND Y = 122 else
"110111011111" when X = 249 AND Y = 122 else
"110111011111" when X = 250 AND Y = 122 else
"110111011111" when X = 251 AND Y = 122 else
"110111011111" when X = 252 AND Y = 122 else
"110111011111" when X = 253 AND Y = 122 else
"110111011111" when X = 254 AND Y = 122 else
"110111011111" when X = 255 AND Y = 122 else
"110111011111" when X = 256 AND Y = 122 else
"110111011111" when X = 257 AND Y = 122 else
"110111011111" when X = 258 AND Y = 122 else
"110111011111" when X = 259 AND Y = 122 else
"110111011111" when X = 260 AND Y = 122 else
"110111011111" when X = 261 AND Y = 122 else
"110111011111" when X = 262 AND Y = 122 else
"110111011111" when X = 263 AND Y = 122 else
"110111011111" when X = 264 AND Y = 122 else
"110111011111" when X = 265 AND Y = 122 else
"110111011111" when X = 266 AND Y = 122 else
"110111011111" when X = 267 AND Y = 122 else
"110111011111" when X = 268 AND Y = 122 else
"110111011111" when X = 269 AND Y = 122 else
"110111011111" when X = 270 AND Y = 122 else
"110111011111" when X = 271 AND Y = 122 else
"110111011111" when X = 272 AND Y = 122 else
"110111011111" when X = 273 AND Y = 122 else
"110111011111" when X = 274 AND Y = 122 else
"110111011111" when X = 275 AND Y = 122 else
"110111011111" when X = 276 AND Y = 122 else
"110111011111" when X = 277 AND Y = 122 else
"110111011111" when X = 278 AND Y = 122 else
"110111011111" when X = 279 AND Y = 122 else
"110111011111" when X = 280 AND Y = 122 else
"110111011111" when X = 281 AND Y = 122 else
"110111011111" when X = 282 AND Y = 122 else
"110111011111" when X = 283 AND Y = 122 else
"110111011111" when X = 284 AND Y = 122 else
"110111011111" when X = 285 AND Y = 122 else
"110111011111" when X = 286 AND Y = 122 else
"110111011111" when X = 287 AND Y = 122 else
"110111011111" when X = 288 AND Y = 122 else
"110111011111" when X = 289 AND Y = 122 else
"110111011111" when X = 290 AND Y = 122 else
"110111011111" when X = 291 AND Y = 122 else
"110111011111" when X = 292 AND Y = 122 else
"110111011111" when X = 293 AND Y = 122 else
"110111011111" when X = 294 AND Y = 122 else
"110111011111" when X = 295 AND Y = 122 else
"110111011111" when X = 296 AND Y = 122 else
"110111011111" when X = 297 AND Y = 122 else
"110111011111" when X = 298 AND Y = 122 else
"110111011111" when X = 299 AND Y = 122 else
"110111011111" when X = 300 AND Y = 122 else
"110111011111" when X = 301 AND Y = 122 else
"110111011111" when X = 302 AND Y = 122 else
"110111011111" when X = 303 AND Y = 122 else
"110111011111" when X = 304 AND Y = 122 else
"110111011111" when X = 305 AND Y = 122 else
"110111011111" when X = 306 AND Y = 122 else
"110111011111" when X = 307 AND Y = 122 else
"110111011111" when X = 308 AND Y = 122 else
"110111011111" when X = 309 AND Y = 122 else
"110111011111" when X = 310 AND Y = 122 else
"110111011111" when X = 311 AND Y = 122 else
"110111011111" when X = 312 AND Y = 122 else
"110111011111" when X = 313 AND Y = 122 else
"110111011111" when X = 314 AND Y = 122 else
"110111011111" when X = 315 AND Y = 122 else
"110111011111" when X = 316 AND Y = 122 else
"110111011111" when X = 317 AND Y = 122 else
"110111011111" when X = 318 AND Y = 122 else
"110111011111" when X = 319 AND Y = 122 else
"110111011111" when X = 320 AND Y = 122 else
"110111011111" when X = 321 AND Y = 122 else
"110111011111" when X = 322 AND Y = 122 else
"110111011111" when X = 323 AND Y = 122 else
"110111011111" when X = 324 AND Y = 122 else
"100010011101" when X = 0 AND Y = 123 else
"100010011101" when X = 1 AND Y = 123 else
"100010011101" when X = 2 AND Y = 123 else
"100010011101" when X = 3 AND Y = 123 else
"100010011101" when X = 4 AND Y = 123 else
"100010011101" when X = 5 AND Y = 123 else
"100010011101" when X = 6 AND Y = 123 else
"100010011101" when X = 7 AND Y = 123 else
"100010011101" when X = 8 AND Y = 123 else
"100010011101" when X = 9 AND Y = 123 else
"100010011101" when X = 10 AND Y = 123 else
"100010011101" when X = 11 AND Y = 123 else
"100010011101" when X = 12 AND Y = 123 else
"100010011101" when X = 13 AND Y = 123 else
"100010011101" when X = 14 AND Y = 123 else
"100010011101" when X = 15 AND Y = 123 else
"100010011101" when X = 16 AND Y = 123 else
"100010011101" when X = 17 AND Y = 123 else
"100010011101" when X = 18 AND Y = 123 else
"100010011101" when X = 19 AND Y = 123 else
"100010011101" when X = 20 AND Y = 123 else
"100010011101" when X = 21 AND Y = 123 else
"100010011101" when X = 22 AND Y = 123 else
"100010011101" when X = 23 AND Y = 123 else
"100010011101" when X = 24 AND Y = 123 else
"100010011101" when X = 25 AND Y = 123 else
"100010011101" when X = 26 AND Y = 123 else
"100010011101" when X = 27 AND Y = 123 else
"100010011101" when X = 28 AND Y = 123 else
"100010011101" when X = 29 AND Y = 123 else
"100010011101" when X = 30 AND Y = 123 else
"100010011101" when X = 31 AND Y = 123 else
"100010011101" when X = 32 AND Y = 123 else
"100010011101" when X = 33 AND Y = 123 else
"100010011101" when X = 34 AND Y = 123 else
"100010011101" when X = 35 AND Y = 123 else
"100010011101" when X = 36 AND Y = 123 else
"100010011101" when X = 37 AND Y = 123 else
"100010011101" when X = 38 AND Y = 123 else
"100010011101" when X = 39 AND Y = 123 else
"110111011111" when X = 40 AND Y = 123 else
"110111011111" when X = 41 AND Y = 123 else
"110111011111" when X = 42 AND Y = 123 else
"110111011111" when X = 43 AND Y = 123 else
"110111011111" when X = 44 AND Y = 123 else
"110111011111" when X = 45 AND Y = 123 else
"110111011111" when X = 46 AND Y = 123 else
"110111011111" when X = 47 AND Y = 123 else
"110111011111" when X = 48 AND Y = 123 else
"110111011111" when X = 49 AND Y = 123 else
"110111011111" when X = 50 AND Y = 123 else
"110111011111" when X = 51 AND Y = 123 else
"110111011111" when X = 52 AND Y = 123 else
"110111011111" when X = 53 AND Y = 123 else
"110111011111" when X = 54 AND Y = 123 else
"110111011111" when X = 55 AND Y = 123 else
"110111011111" when X = 56 AND Y = 123 else
"110111011111" when X = 57 AND Y = 123 else
"110111011111" when X = 58 AND Y = 123 else
"110111011111" when X = 59 AND Y = 123 else
"110111011111" when X = 60 AND Y = 123 else
"110111011111" when X = 61 AND Y = 123 else
"110111011111" when X = 62 AND Y = 123 else
"110111011111" when X = 63 AND Y = 123 else
"110111011111" when X = 64 AND Y = 123 else
"110111011111" when X = 65 AND Y = 123 else
"110111011111" when X = 66 AND Y = 123 else
"110111011111" when X = 67 AND Y = 123 else
"110111011111" when X = 68 AND Y = 123 else
"110111011111" when X = 69 AND Y = 123 else
"110111011111" when X = 70 AND Y = 123 else
"110111011111" when X = 71 AND Y = 123 else
"110111011111" when X = 72 AND Y = 123 else
"110111011111" when X = 73 AND Y = 123 else
"110111011111" when X = 74 AND Y = 123 else
"110111011111" when X = 75 AND Y = 123 else
"110111011111" when X = 76 AND Y = 123 else
"110111011111" when X = 77 AND Y = 123 else
"110111011111" when X = 78 AND Y = 123 else
"110111011111" when X = 79 AND Y = 123 else
"110111011111" when X = 80 AND Y = 123 else
"110111011111" when X = 81 AND Y = 123 else
"110111011111" when X = 82 AND Y = 123 else
"110111011111" when X = 83 AND Y = 123 else
"110111011111" when X = 84 AND Y = 123 else
"110111011111" when X = 85 AND Y = 123 else
"110111011111" when X = 86 AND Y = 123 else
"110111011111" when X = 87 AND Y = 123 else
"110111011111" when X = 88 AND Y = 123 else
"110111011111" when X = 89 AND Y = 123 else
"110111011111" when X = 90 AND Y = 123 else
"110111011111" when X = 91 AND Y = 123 else
"110111011111" when X = 92 AND Y = 123 else
"110111011111" when X = 93 AND Y = 123 else
"110111011111" when X = 94 AND Y = 123 else
"110111011111" when X = 95 AND Y = 123 else
"110111011111" when X = 96 AND Y = 123 else
"110111011111" when X = 97 AND Y = 123 else
"110111011111" when X = 98 AND Y = 123 else
"110111011111" when X = 99 AND Y = 123 else
"110111011111" when X = 100 AND Y = 123 else
"110111011111" when X = 101 AND Y = 123 else
"110111011111" when X = 102 AND Y = 123 else
"110111011111" when X = 103 AND Y = 123 else
"110111011111" when X = 104 AND Y = 123 else
"110111011111" when X = 105 AND Y = 123 else
"110111011111" when X = 106 AND Y = 123 else
"110111011111" when X = 107 AND Y = 123 else
"110111011111" when X = 108 AND Y = 123 else
"110111011111" when X = 109 AND Y = 123 else
"110111011111" when X = 110 AND Y = 123 else
"110111011111" when X = 111 AND Y = 123 else
"110111011111" when X = 112 AND Y = 123 else
"110111011111" when X = 113 AND Y = 123 else
"110111011111" when X = 114 AND Y = 123 else
"110111011111" when X = 115 AND Y = 123 else
"110111011111" when X = 116 AND Y = 123 else
"110111011111" when X = 117 AND Y = 123 else
"110111011111" when X = 118 AND Y = 123 else
"110111011111" when X = 119 AND Y = 123 else
"110111011111" when X = 120 AND Y = 123 else
"110111011111" when X = 121 AND Y = 123 else
"110111011111" when X = 122 AND Y = 123 else
"110111011111" when X = 123 AND Y = 123 else
"110111011111" when X = 124 AND Y = 123 else
"110111011111" when X = 125 AND Y = 123 else
"110111011111" when X = 126 AND Y = 123 else
"110111011111" when X = 127 AND Y = 123 else
"110111011111" when X = 128 AND Y = 123 else
"110111011111" when X = 129 AND Y = 123 else
"110111011111" when X = 130 AND Y = 123 else
"110111011111" when X = 131 AND Y = 123 else
"110111011111" when X = 132 AND Y = 123 else
"110111011111" when X = 133 AND Y = 123 else
"110111011111" when X = 134 AND Y = 123 else
"110111011111" when X = 135 AND Y = 123 else
"110111011111" when X = 136 AND Y = 123 else
"110111011111" when X = 137 AND Y = 123 else
"110111011111" when X = 138 AND Y = 123 else
"110111011111" when X = 139 AND Y = 123 else
"110111011111" when X = 140 AND Y = 123 else
"110111011111" when X = 141 AND Y = 123 else
"110111011111" when X = 142 AND Y = 123 else
"110111011111" when X = 143 AND Y = 123 else
"110111011111" when X = 144 AND Y = 123 else
"110111011111" when X = 145 AND Y = 123 else
"110111011111" when X = 146 AND Y = 123 else
"110111011111" when X = 147 AND Y = 123 else
"110111011111" when X = 148 AND Y = 123 else
"110111011111" when X = 149 AND Y = 123 else
"110111011111" when X = 150 AND Y = 123 else
"110111011111" when X = 151 AND Y = 123 else
"110111011111" when X = 152 AND Y = 123 else
"110111011111" when X = 153 AND Y = 123 else
"110111011111" when X = 154 AND Y = 123 else
"110111011111" when X = 155 AND Y = 123 else
"110111011111" when X = 156 AND Y = 123 else
"110111011111" when X = 157 AND Y = 123 else
"110111011111" when X = 158 AND Y = 123 else
"110111011111" when X = 159 AND Y = 123 else
"110111011111" when X = 160 AND Y = 123 else
"110111011111" when X = 161 AND Y = 123 else
"110111011111" when X = 162 AND Y = 123 else
"110111011111" when X = 163 AND Y = 123 else
"110111011111" when X = 164 AND Y = 123 else
"111111111111" when X = 165 AND Y = 123 else
"111111111111" when X = 166 AND Y = 123 else
"111111111111" when X = 167 AND Y = 123 else
"111111111111" when X = 168 AND Y = 123 else
"111111111111" when X = 169 AND Y = 123 else
"111111111111" when X = 170 AND Y = 123 else
"111111111111" when X = 171 AND Y = 123 else
"111111111111" when X = 172 AND Y = 123 else
"111111111111" when X = 173 AND Y = 123 else
"111111111111" when X = 174 AND Y = 123 else
"111111111111" when X = 175 AND Y = 123 else
"111111111111" when X = 176 AND Y = 123 else
"111111111111" when X = 177 AND Y = 123 else
"111111111111" when X = 178 AND Y = 123 else
"111111111111" when X = 179 AND Y = 123 else
"111111111111" when X = 180 AND Y = 123 else
"111111111111" when X = 181 AND Y = 123 else
"111111111111" when X = 182 AND Y = 123 else
"111111111111" when X = 183 AND Y = 123 else
"111111111111" when X = 184 AND Y = 123 else
"111111111111" when X = 185 AND Y = 123 else
"111111111111" when X = 186 AND Y = 123 else
"111111111111" when X = 187 AND Y = 123 else
"111111111111" when X = 188 AND Y = 123 else
"111111111111" when X = 189 AND Y = 123 else
"110111011111" when X = 190 AND Y = 123 else
"110111011111" when X = 191 AND Y = 123 else
"110111011111" when X = 192 AND Y = 123 else
"110111011111" when X = 193 AND Y = 123 else
"110111011111" when X = 194 AND Y = 123 else
"110111011111" when X = 195 AND Y = 123 else
"110111011111" when X = 196 AND Y = 123 else
"110111011111" when X = 197 AND Y = 123 else
"110111011111" when X = 198 AND Y = 123 else
"110111011111" when X = 199 AND Y = 123 else
"110111011111" when X = 200 AND Y = 123 else
"110111011111" when X = 201 AND Y = 123 else
"110111011111" when X = 202 AND Y = 123 else
"110111011111" when X = 203 AND Y = 123 else
"110111011111" when X = 204 AND Y = 123 else
"110111011111" when X = 205 AND Y = 123 else
"110111011111" when X = 206 AND Y = 123 else
"110111011111" when X = 207 AND Y = 123 else
"110111011111" when X = 208 AND Y = 123 else
"110111011111" when X = 209 AND Y = 123 else
"110111011111" when X = 210 AND Y = 123 else
"110111011111" when X = 211 AND Y = 123 else
"110111011111" when X = 212 AND Y = 123 else
"110111011111" when X = 213 AND Y = 123 else
"110111011111" when X = 214 AND Y = 123 else
"110111011111" when X = 215 AND Y = 123 else
"110111011111" when X = 216 AND Y = 123 else
"110111011111" when X = 217 AND Y = 123 else
"110111011111" when X = 218 AND Y = 123 else
"110111011111" when X = 219 AND Y = 123 else
"110111011111" when X = 220 AND Y = 123 else
"110111011111" when X = 221 AND Y = 123 else
"110111011111" when X = 222 AND Y = 123 else
"110111011111" when X = 223 AND Y = 123 else
"110111011111" when X = 224 AND Y = 123 else
"110111011111" when X = 225 AND Y = 123 else
"110111011111" when X = 226 AND Y = 123 else
"110111011111" when X = 227 AND Y = 123 else
"110111011111" when X = 228 AND Y = 123 else
"110111011111" when X = 229 AND Y = 123 else
"110111011111" when X = 230 AND Y = 123 else
"110111011111" when X = 231 AND Y = 123 else
"110111011111" when X = 232 AND Y = 123 else
"110111011111" when X = 233 AND Y = 123 else
"110111011111" when X = 234 AND Y = 123 else
"110111011111" when X = 235 AND Y = 123 else
"110111011111" when X = 236 AND Y = 123 else
"110111011111" when X = 237 AND Y = 123 else
"110111011111" when X = 238 AND Y = 123 else
"110111011111" when X = 239 AND Y = 123 else
"110111011111" when X = 240 AND Y = 123 else
"110111011111" when X = 241 AND Y = 123 else
"110111011111" when X = 242 AND Y = 123 else
"110111011111" when X = 243 AND Y = 123 else
"110111011111" when X = 244 AND Y = 123 else
"110111011111" when X = 245 AND Y = 123 else
"110111011111" when X = 246 AND Y = 123 else
"110111011111" when X = 247 AND Y = 123 else
"110111011111" when X = 248 AND Y = 123 else
"110111011111" when X = 249 AND Y = 123 else
"110111011111" when X = 250 AND Y = 123 else
"110111011111" when X = 251 AND Y = 123 else
"110111011111" when X = 252 AND Y = 123 else
"110111011111" when X = 253 AND Y = 123 else
"110111011111" when X = 254 AND Y = 123 else
"110111011111" when X = 255 AND Y = 123 else
"110111011111" when X = 256 AND Y = 123 else
"110111011111" when X = 257 AND Y = 123 else
"110111011111" when X = 258 AND Y = 123 else
"110111011111" when X = 259 AND Y = 123 else
"110111011111" when X = 260 AND Y = 123 else
"110111011111" when X = 261 AND Y = 123 else
"110111011111" when X = 262 AND Y = 123 else
"110111011111" when X = 263 AND Y = 123 else
"110111011111" when X = 264 AND Y = 123 else
"110111011111" when X = 265 AND Y = 123 else
"110111011111" when X = 266 AND Y = 123 else
"110111011111" when X = 267 AND Y = 123 else
"110111011111" when X = 268 AND Y = 123 else
"110111011111" when X = 269 AND Y = 123 else
"110111011111" when X = 270 AND Y = 123 else
"110111011111" when X = 271 AND Y = 123 else
"110111011111" when X = 272 AND Y = 123 else
"110111011111" when X = 273 AND Y = 123 else
"110111011111" when X = 274 AND Y = 123 else
"110111011111" when X = 275 AND Y = 123 else
"110111011111" when X = 276 AND Y = 123 else
"110111011111" when X = 277 AND Y = 123 else
"110111011111" when X = 278 AND Y = 123 else
"110111011111" when X = 279 AND Y = 123 else
"110111011111" when X = 280 AND Y = 123 else
"110111011111" when X = 281 AND Y = 123 else
"110111011111" when X = 282 AND Y = 123 else
"110111011111" when X = 283 AND Y = 123 else
"110111011111" when X = 284 AND Y = 123 else
"110111011111" when X = 285 AND Y = 123 else
"110111011111" when X = 286 AND Y = 123 else
"110111011111" when X = 287 AND Y = 123 else
"110111011111" when X = 288 AND Y = 123 else
"110111011111" when X = 289 AND Y = 123 else
"110111011111" when X = 290 AND Y = 123 else
"110111011111" when X = 291 AND Y = 123 else
"110111011111" when X = 292 AND Y = 123 else
"110111011111" when X = 293 AND Y = 123 else
"110111011111" when X = 294 AND Y = 123 else
"110111011111" when X = 295 AND Y = 123 else
"110111011111" when X = 296 AND Y = 123 else
"110111011111" when X = 297 AND Y = 123 else
"110111011111" when X = 298 AND Y = 123 else
"110111011111" when X = 299 AND Y = 123 else
"110111011111" when X = 300 AND Y = 123 else
"110111011111" when X = 301 AND Y = 123 else
"110111011111" when X = 302 AND Y = 123 else
"110111011111" when X = 303 AND Y = 123 else
"110111011111" when X = 304 AND Y = 123 else
"110111011111" when X = 305 AND Y = 123 else
"110111011111" when X = 306 AND Y = 123 else
"110111011111" when X = 307 AND Y = 123 else
"110111011111" when X = 308 AND Y = 123 else
"110111011111" when X = 309 AND Y = 123 else
"110111011111" when X = 310 AND Y = 123 else
"110111011111" when X = 311 AND Y = 123 else
"110111011111" when X = 312 AND Y = 123 else
"110111011111" when X = 313 AND Y = 123 else
"110111011111" when X = 314 AND Y = 123 else
"110111011111" when X = 315 AND Y = 123 else
"110111011111" when X = 316 AND Y = 123 else
"110111011111" when X = 317 AND Y = 123 else
"110111011111" when X = 318 AND Y = 123 else
"110111011111" when X = 319 AND Y = 123 else
"110111011111" when X = 320 AND Y = 123 else
"110111011111" when X = 321 AND Y = 123 else
"110111011111" when X = 322 AND Y = 123 else
"110111011111" when X = 323 AND Y = 123 else
"110111011111" when X = 324 AND Y = 123 else
"100010011101" when X = 0 AND Y = 124 else
"100010011101" when X = 1 AND Y = 124 else
"100010011101" when X = 2 AND Y = 124 else
"100010011101" when X = 3 AND Y = 124 else
"100010011101" when X = 4 AND Y = 124 else
"100010011101" when X = 5 AND Y = 124 else
"100010011101" when X = 6 AND Y = 124 else
"100010011101" when X = 7 AND Y = 124 else
"100010011101" when X = 8 AND Y = 124 else
"100010011101" when X = 9 AND Y = 124 else
"100010011101" when X = 10 AND Y = 124 else
"100010011101" when X = 11 AND Y = 124 else
"100010011101" when X = 12 AND Y = 124 else
"100010011101" when X = 13 AND Y = 124 else
"100010011101" when X = 14 AND Y = 124 else
"100010011101" when X = 15 AND Y = 124 else
"100010011101" when X = 16 AND Y = 124 else
"100010011101" when X = 17 AND Y = 124 else
"100010011101" when X = 18 AND Y = 124 else
"100010011101" when X = 19 AND Y = 124 else
"100010011101" when X = 20 AND Y = 124 else
"100010011101" when X = 21 AND Y = 124 else
"100010011101" when X = 22 AND Y = 124 else
"100010011101" when X = 23 AND Y = 124 else
"100010011101" when X = 24 AND Y = 124 else
"100010011101" when X = 25 AND Y = 124 else
"100010011101" when X = 26 AND Y = 124 else
"100010011101" when X = 27 AND Y = 124 else
"100010011101" when X = 28 AND Y = 124 else
"100010011101" when X = 29 AND Y = 124 else
"100010011101" when X = 30 AND Y = 124 else
"100010011101" when X = 31 AND Y = 124 else
"100010011101" when X = 32 AND Y = 124 else
"100010011101" when X = 33 AND Y = 124 else
"100010011101" when X = 34 AND Y = 124 else
"100010011101" when X = 35 AND Y = 124 else
"100010011101" when X = 36 AND Y = 124 else
"100010011101" when X = 37 AND Y = 124 else
"100010011101" when X = 38 AND Y = 124 else
"100010011101" when X = 39 AND Y = 124 else
"110111011111" when X = 40 AND Y = 124 else
"110111011111" when X = 41 AND Y = 124 else
"110111011111" when X = 42 AND Y = 124 else
"110111011111" when X = 43 AND Y = 124 else
"110111011111" when X = 44 AND Y = 124 else
"110111011111" when X = 45 AND Y = 124 else
"110111011111" when X = 46 AND Y = 124 else
"110111011111" when X = 47 AND Y = 124 else
"110111011111" when X = 48 AND Y = 124 else
"110111011111" when X = 49 AND Y = 124 else
"110111011111" when X = 50 AND Y = 124 else
"110111011111" when X = 51 AND Y = 124 else
"110111011111" when X = 52 AND Y = 124 else
"110111011111" when X = 53 AND Y = 124 else
"110111011111" when X = 54 AND Y = 124 else
"110111011111" when X = 55 AND Y = 124 else
"110111011111" when X = 56 AND Y = 124 else
"110111011111" when X = 57 AND Y = 124 else
"110111011111" when X = 58 AND Y = 124 else
"110111011111" when X = 59 AND Y = 124 else
"110111011111" when X = 60 AND Y = 124 else
"110111011111" when X = 61 AND Y = 124 else
"110111011111" when X = 62 AND Y = 124 else
"110111011111" when X = 63 AND Y = 124 else
"110111011111" when X = 64 AND Y = 124 else
"110111011111" when X = 65 AND Y = 124 else
"110111011111" when X = 66 AND Y = 124 else
"110111011111" when X = 67 AND Y = 124 else
"110111011111" when X = 68 AND Y = 124 else
"110111011111" when X = 69 AND Y = 124 else
"110111011111" when X = 70 AND Y = 124 else
"110111011111" when X = 71 AND Y = 124 else
"110111011111" when X = 72 AND Y = 124 else
"110111011111" when X = 73 AND Y = 124 else
"110111011111" when X = 74 AND Y = 124 else
"110111011111" when X = 75 AND Y = 124 else
"110111011111" when X = 76 AND Y = 124 else
"110111011111" when X = 77 AND Y = 124 else
"110111011111" when X = 78 AND Y = 124 else
"110111011111" when X = 79 AND Y = 124 else
"110111011111" when X = 80 AND Y = 124 else
"110111011111" when X = 81 AND Y = 124 else
"110111011111" when X = 82 AND Y = 124 else
"110111011111" when X = 83 AND Y = 124 else
"110111011111" when X = 84 AND Y = 124 else
"110111011111" when X = 85 AND Y = 124 else
"110111011111" when X = 86 AND Y = 124 else
"110111011111" when X = 87 AND Y = 124 else
"110111011111" when X = 88 AND Y = 124 else
"110111011111" when X = 89 AND Y = 124 else
"110111011111" when X = 90 AND Y = 124 else
"110111011111" when X = 91 AND Y = 124 else
"110111011111" when X = 92 AND Y = 124 else
"110111011111" when X = 93 AND Y = 124 else
"110111011111" when X = 94 AND Y = 124 else
"110111011111" when X = 95 AND Y = 124 else
"110111011111" when X = 96 AND Y = 124 else
"110111011111" when X = 97 AND Y = 124 else
"110111011111" when X = 98 AND Y = 124 else
"110111011111" when X = 99 AND Y = 124 else
"110111011111" when X = 100 AND Y = 124 else
"110111011111" when X = 101 AND Y = 124 else
"110111011111" when X = 102 AND Y = 124 else
"110111011111" when X = 103 AND Y = 124 else
"110111011111" when X = 104 AND Y = 124 else
"110111011111" when X = 105 AND Y = 124 else
"110111011111" when X = 106 AND Y = 124 else
"110111011111" when X = 107 AND Y = 124 else
"110111011111" when X = 108 AND Y = 124 else
"110111011111" when X = 109 AND Y = 124 else
"110111011111" when X = 110 AND Y = 124 else
"110111011111" when X = 111 AND Y = 124 else
"110111011111" when X = 112 AND Y = 124 else
"110111011111" when X = 113 AND Y = 124 else
"110111011111" when X = 114 AND Y = 124 else
"110111011111" when X = 115 AND Y = 124 else
"110111011111" when X = 116 AND Y = 124 else
"110111011111" when X = 117 AND Y = 124 else
"110111011111" when X = 118 AND Y = 124 else
"110111011111" when X = 119 AND Y = 124 else
"110111011111" when X = 120 AND Y = 124 else
"110111011111" when X = 121 AND Y = 124 else
"110111011111" when X = 122 AND Y = 124 else
"110111011111" when X = 123 AND Y = 124 else
"110111011111" when X = 124 AND Y = 124 else
"110111011111" when X = 125 AND Y = 124 else
"110111011111" when X = 126 AND Y = 124 else
"110111011111" when X = 127 AND Y = 124 else
"110111011111" when X = 128 AND Y = 124 else
"110111011111" when X = 129 AND Y = 124 else
"110111011111" when X = 130 AND Y = 124 else
"110111011111" when X = 131 AND Y = 124 else
"110111011111" when X = 132 AND Y = 124 else
"110111011111" when X = 133 AND Y = 124 else
"110111011111" when X = 134 AND Y = 124 else
"110111011111" when X = 135 AND Y = 124 else
"110111011111" when X = 136 AND Y = 124 else
"110111011111" when X = 137 AND Y = 124 else
"110111011111" when X = 138 AND Y = 124 else
"110111011111" when X = 139 AND Y = 124 else
"110111011111" when X = 140 AND Y = 124 else
"110111011111" when X = 141 AND Y = 124 else
"110111011111" when X = 142 AND Y = 124 else
"110111011111" when X = 143 AND Y = 124 else
"110111011111" when X = 144 AND Y = 124 else
"110111011111" when X = 145 AND Y = 124 else
"110111011111" when X = 146 AND Y = 124 else
"110111011111" when X = 147 AND Y = 124 else
"110111011111" when X = 148 AND Y = 124 else
"110111011111" when X = 149 AND Y = 124 else
"110111011111" when X = 150 AND Y = 124 else
"110111011111" when X = 151 AND Y = 124 else
"110111011111" when X = 152 AND Y = 124 else
"110111011111" when X = 153 AND Y = 124 else
"110111011111" when X = 154 AND Y = 124 else
"110111011111" when X = 155 AND Y = 124 else
"110111011111" when X = 156 AND Y = 124 else
"110111011111" when X = 157 AND Y = 124 else
"110111011111" when X = 158 AND Y = 124 else
"110111011111" when X = 159 AND Y = 124 else
"110111011111" when X = 160 AND Y = 124 else
"110111011111" when X = 161 AND Y = 124 else
"110111011111" when X = 162 AND Y = 124 else
"110111011111" when X = 163 AND Y = 124 else
"110111011111" when X = 164 AND Y = 124 else
"111111111111" when X = 165 AND Y = 124 else
"111111111111" when X = 166 AND Y = 124 else
"111111111111" when X = 167 AND Y = 124 else
"111111111111" when X = 168 AND Y = 124 else
"111111111111" when X = 169 AND Y = 124 else
"111111111111" when X = 170 AND Y = 124 else
"111111111111" when X = 171 AND Y = 124 else
"111111111111" when X = 172 AND Y = 124 else
"111111111111" when X = 173 AND Y = 124 else
"111111111111" when X = 174 AND Y = 124 else
"111111111111" when X = 175 AND Y = 124 else
"111111111111" when X = 176 AND Y = 124 else
"111111111111" when X = 177 AND Y = 124 else
"111111111111" when X = 178 AND Y = 124 else
"111111111111" when X = 179 AND Y = 124 else
"111111111111" when X = 180 AND Y = 124 else
"111111111111" when X = 181 AND Y = 124 else
"111111111111" when X = 182 AND Y = 124 else
"111111111111" when X = 183 AND Y = 124 else
"111111111111" when X = 184 AND Y = 124 else
"111111111111" when X = 185 AND Y = 124 else
"111111111111" when X = 186 AND Y = 124 else
"111111111111" when X = 187 AND Y = 124 else
"111111111111" when X = 188 AND Y = 124 else
"111111111111" when X = 189 AND Y = 124 else
"110111011111" when X = 190 AND Y = 124 else
"110111011111" when X = 191 AND Y = 124 else
"110111011111" when X = 192 AND Y = 124 else
"110111011111" when X = 193 AND Y = 124 else
"110111011111" when X = 194 AND Y = 124 else
"110111011111" when X = 195 AND Y = 124 else
"110111011111" when X = 196 AND Y = 124 else
"110111011111" when X = 197 AND Y = 124 else
"110111011111" when X = 198 AND Y = 124 else
"110111011111" when X = 199 AND Y = 124 else
"110111011111" when X = 200 AND Y = 124 else
"110111011111" when X = 201 AND Y = 124 else
"110111011111" when X = 202 AND Y = 124 else
"110111011111" when X = 203 AND Y = 124 else
"110111011111" when X = 204 AND Y = 124 else
"110111011111" when X = 205 AND Y = 124 else
"110111011111" when X = 206 AND Y = 124 else
"110111011111" when X = 207 AND Y = 124 else
"110111011111" when X = 208 AND Y = 124 else
"110111011111" when X = 209 AND Y = 124 else
"110111011111" when X = 210 AND Y = 124 else
"110111011111" when X = 211 AND Y = 124 else
"110111011111" when X = 212 AND Y = 124 else
"110111011111" when X = 213 AND Y = 124 else
"110111011111" when X = 214 AND Y = 124 else
"110111011111" when X = 215 AND Y = 124 else
"110111011111" when X = 216 AND Y = 124 else
"110111011111" when X = 217 AND Y = 124 else
"110111011111" when X = 218 AND Y = 124 else
"110111011111" when X = 219 AND Y = 124 else
"110111011111" when X = 220 AND Y = 124 else
"110111011111" when X = 221 AND Y = 124 else
"110111011111" when X = 222 AND Y = 124 else
"110111011111" when X = 223 AND Y = 124 else
"110111011111" when X = 224 AND Y = 124 else
"110111011111" when X = 225 AND Y = 124 else
"110111011111" when X = 226 AND Y = 124 else
"110111011111" when X = 227 AND Y = 124 else
"110111011111" when X = 228 AND Y = 124 else
"110111011111" when X = 229 AND Y = 124 else
"110111011111" when X = 230 AND Y = 124 else
"110111011111" when X = 231 AND Y = 124 else
"110111011111" when X = 232 AND Y = 124 else
"110111011111" when X = 233 AND Y = 124 else
"110111011111" when X = 234 AND Y = 124 else
"110111011111" when X = 235 AND Y = 124 else
"110111011111" when X = 236 AND Y = 124 else
"110111011111" when X = 237 AND Y = 124 else
"110111011111" when X = 238 AND Y = 124 else
"110111011111" when X = 239 AND Y = 124 else
"110111011111" when X = 240 AND Y = 124 else
"110111011111" when X = 241 AND Y = 124 else
"110111011111" when X = 242 AND Y = 124 else
"110111011111" when X = 243 AND Y = 124 else
"110111011111" when X = 244 AND Y = 124 else
"110111011111" when X = 245 AND Y = 124 else
"110111011111" when X = 246 AND Y = 124 else
"110111011111" when X = 247 AND Y = 124 else
"110111011111" when X = 248 AND Y = 124 else
"110111011111" when X = 249 AND Y = 124 else
"110111011111" when X = 250 AND Y = 124 else
"110111011111" when X = 251 AND Y = 124 else
"110111011111" when X = 252 AND Y = 124 else
"110111011111" when X = 253 AND Y = 124 else
"110111011111" when X = 254 AND Y = 124 else
"110111011111" when X = 255 AND Y = 124 else
"110111011111" when X = 256 AND Y = 124 else
"110111011111" when X = 257 AND Y = 124 else
"110111011111" when X = 258 AND Y = 124 else
"110111011111" when X = 259 AND Y = 124 else
"110111011111" when X = 260 AND Y = 124 else
"110111011111" when X = 261 AND Y = 124 else
"110111011111" when X = 262 AND Y = 124 else
"110111011111" when X = 263 AND Y = 124 else
"110111011111" when X = 264 AND Y = 124 else
"110111011111" when X = 265 AND Y = 124 else
"110111011111" when X = 266 AND Y = 124 else
"110111011111" when X = 267 AND Y = 124 else
"110111011111" when X = 268 AND Y = 124 else
"110111011111" when X = 269 AND Y = 124 else
"110111011111" when X = 270 AND Y = 124 else
"110111011111" when X = 271 AND Y = 124 else
"110111011111" when X = 272 AND Y = 124 else
"110111011111" when X = 273 AND Y = 124 else
"110111011111" when X = 274 AND Y = 124 else
"110111011111" when X = 275 AND Y = 124 else
"110111011111" when X = 276 AND Y = 124 else
"110111011111" when X = 277 AND Y = 124 else
"110111011111" when X = 278 AND Y = 124 else
"110111011111" when X = 279 AND Y = 124 else
"110111011111" when X = 280 AND Y = 124 else
"110111011111" when X = 281 AND Y = 124 else
"110111011111" when X = 282 AND Y = 124 else
"110111011111" when X = 283 AND Y = 124 else
"110111011111" when X = 284 AND Y = 124 else
"110111011111" when X = 285 AND Y = 124 else
"110111011111" when X = 286 AND Y = 124 else
"110111011111" when X = 287 AND Y = 124 else
"110111011111" when X = 288 AND Y = 124 else
"110111011111" when X = 289 AND Y = 124 else
"110111011111" when X = 290 AND Y = 124 else
"110111011111" when X = 291 AND Y = 124 else
"110111011111" when X = 292 AND Y = 124 else
"110111011111" when X = 293 AND Y = 124 else
"110111011111" when X = 294 AND Y = 124 else
"110111011111" when X = 295 AND Y = 124 else
"110111011111" when X = 296 AND Y = 124 else
"110111011111" when X = 297 AND Y = 124 else
"110111011111" when X = 298 AND Y = 124 else
"110111011111" when X = 299 AND Y = 124 else
"110111011111" when X = 300 AND Y = 124 else
"110111011111" when X = 301 AND Y = 124 else
"110111011111" when X = 302 AND Y = 124 else
"110111011111" when X = 303 AND Y = 124 else
"110111011111" when X = 304 AND Y = 124 else
"110111011111" when X = 305 AND Y = 124 else
"110111011111" when X = 306 AND Y = 124 else
"110111011111" when X = 307 AND Y = 124 else
"110111011111" when X = 308 AND Y = 124 else
"110111011111" when X = 309 AND Y = 124 else
"110111011111" when X = 310 AND Y = 124 else
"110111011111" when X = 311 AND Y = 124 else
"110111011111" when X = 312 AND Y = 124 else
"110111011111" when X = 313 AND Y = 124 else
"110111011111" when X = 314 AND Y = 124 else
"110111011111" when X = 315 AND Y = 124 else
"110111011111" when X = 316 AND Y = 124 else
"110111011111" when X = 317 AND Y = 124 else
"110111011111" when X = 318 AND Y = 124 else
"110111011111" when X = 319 AND Y = 124 else
"110111011111" when X = 320 AND Y = 124 else
"110111011111" when X = 321 AND Y = 124 else
"110111011111" when X = 322 AND Y = 124 else
"110111011111" when X = 323 AND Y = 124 else
"110111011111" when X = 324 AND Y = 124 else
"100010011101" when X = 0 AND Y = 125 else
"100010011101" when X = 1 AND Y = 125 else
"100010011101" when X = 2 AND Y = 125 else
"100010011101" when X = 3 AND Y = 125 else
"100010011101" when X = 4 AND Y = 125 else
"100010011101" when X = 5 AND Y = 125 else
"100010011101" when X = 6 AND Y = 125 else
"100010011101" when X = 7 AND Y = 125 else
"100010011101" when X = 8 AND Y = 125 else
"100010011101" when X = 9 AND Y = 125 else
"100010011101" when X = 10 AND Y = 125 else
"100010011101" when X = 11 AND Y = 125 else
"100010011101" when X = 12 AND Y = 125 else
"100010011101" when X = 13 AND Y = 125 else
"100010011101" when X = 14 AND Y = 125 else
"100010011101" when X = 15 AND Y = 125 else
"100010011101" when X = 16 AND Y = 125 else
"100010011101" when X = 17 AND Y = 125 else
"100010011101" when X = 18 AND Y = 125 else
"100010011101" when X = 19 AND Y = 125 else
"100010011101" when X = 20 AND Y = 125 else
"100010011101" when X = 21 AND Y = 125 else
"100010011101" when X = 22 AND Y = 125 else
"100010011101" when X = 23 AND Y = 125 else
"100010011101" when X = 24 AND Y = 125 else
"100010011101" when X = 25 AND Y = 125 else
"100010011101" when X = 26 AND Y = 125 else
"100010011101" when X = 27 AND Y = 125 else
"100010011101" when X = 28 AND Y = 125 else
"100010011101" when X = 29 AND Y = 125 else
"100010011101" when X = 30 AND Y = 125 else
"100010011101" when X = 31 AND Y = 125 else
"100010011101" when X = 32 AND Y = 125 else
"100010011101" when X = 33 AND Y = 125 else
"100010011101" when X = 34 AND Y = 125 else
"100010011101" when X = 35 AND Y = 125 else
"100010011101" when X = 36 AND Y = 125 else
"100010011101" when X = 37 AND Y = 125 else
"100010011101" when X = 38 AND Y = 125 else
"100010011101" when X = 39 AND Y = 125 else
"100010011101" when X = 40 AND Y = 125 else
"100010011101" when X = 41 AND Y = 125 else
"100010011101" when X = 42 AND Y = 125 else
"100010011101" when X = 43 AND Y = 125 else
"100010011101" when X = 44 AND Y = 125 else
"100010011101" when X = 45 AND Y = 125 else
"100010011101" when X = 46 AND Y = 125 else
"100010011101" when X = 47 AND Y = 125 else
"100010011101" when X = 48 AND Y = 125 else
"100010011101" when X = 49 AND Y = 125 else
"100010011101" when X = 50 AND Y = 125 else
"100010011101" when X = 51 AND Y = 125 else
"100010011101" when X = 52 AND Y = 125 else
"100010011101" when X = 53 AND Y = 125 else
"100010011101" when X = 54 AND Y = 125 else
"100010011101" when X = 55 AND Y = 125 else
"100010011101" when X = 56 AND Y = 125 else
"100010011101" when X = 57 AND Y = 125 else
"100010011101" when X = 58 AND Y = 125 else
"100010011101" when X = 59 AND Y = 125 else
"100010011101" when X = 60 AND Y = 125 else
"100010011101" when X = 61 AND Y = 125 else
"100010011101" when X = 62 AND Y = 125 else
"100010011101" when X = 63 AND Y = 125 else
"100010011101" when X = 64 AND Y = 125 else
"100010011101" when X = 65 AND Y = 125 else
"100010011101" when X = 66 AND Y = 125 else
"100010011101" when X = 67 AND Y = 125 else
"100010011101" when X = 68 AND Y = 125 else
"100010011101" when X = 69 AND Y = 125 else
"100010011101" when X = 70 AND Y = 125 else
"100010011101" when X = 71 AND Y = 125 else
"100010011101" when X = 72 AND Y = 125 else
"100010011101" when X = 73 AND Y = 125 else
"100010011101" when X = 74 AND Y = 125 else
"100010011101" when X = 75 AND Y = 125 else
"100010011101" when X = 76 AND Y = 125 else
"100010011101" when X = 77 AND Y = 125 else
"100010011101" when X = 78 AND Y = 125 else
"100010011101" when X = 79 AND Y = 125 else
"100010011101" when X = 80 AND Y = 125 else
"100010011101" when X = 81 AND Y = 125 else
"100010011101" when X = 82 AND Y = 125 else
"100010011101" when X = 83 AND Y = 125 else
"100010011101" when X = 84 AND Y = 125 else
"100010011101" when X = 85 AND Y = 125 else
"100010011101" when X = 86 AND Y = 125 else
"100010011101" when X = 87 AND Y = 125 else
"100010011101" when X = 88 AND Y = 125 else
"100010011101" when X = 89 AND Y = 125 else
"100010011101" when X = 90 AND Y = 125 else
"100010011101" when X = 91 AND Y = 125 else
"100010011101" when X = 92 AND Y = 125 else
"100010011101" when X = 93 AND Y = 125 else
"100010011101" when X = 94 AND Y = 125 else
"100010011101" when X = 95 AND Y = 125 else
"100010011101" when X = 96 AND Y = 125 else
"100010011101" when X = 97 AND Y = 125 else
"100010011101" when X = 98 AND Y = 125 else
"100010011101" when X = 99 AND Y = 125 else
"100010011101" when X = 100 AND Y = 125 else
"100010011101" when X = 101 AND Y = 125 else
"100010011101" when X = 102 AND Y = 125 else
"100010011101" when X = 103 AND Y = 125 else
"100010011101" when X = 104 AND Y = 125 else
"100010011101" when X = 105 AND Y = 125 else
"100010011101" when X = 106 AND Y = 125 else
"100010011101" when X = 107 AND Y = 125 else
"100010011101" when X = 108 AND Y = 125 else
"100010011101" when X = 109 AND Y = 125 else
"110111011111" when X = 110 AND Y = 125 else
"110111011111" when X = 111 AND Y = 125 else
"110111011111" when X = 112 AND Y = 125 else
"110111011111" when X = 113 AND Y = 125 else
"110111011111" when X = 114 AND Y = 125 else
"110111011111" when X = 115 AND Y = 125 else
"110111011111" when X = 116 AND Y = 125 else
"110111011111" when X = 117 AND Y = 125 else
"110111011111" when X = 118 AND Y = 125 else
"110111011111" when X = 119 AND Y = 125 else
"110111011111" when X = 120 AND Y = 125 else
"110111011111" when X = 121 AND Y = 125 else
"110111011111" when X = 122 AND Y = 125 else
"110111011111" when X = 123 AND Y = 125 else
"110111011111" when X = 124 AND Y = 125 else
"110111011111" when X = 125 AND Y = 125 else
"110111011111" when X = 126 AND Y = 125 else
"110111011111" when X = 127 AND Y = 125 else
"110111011111" when X = 128 AND Y = 125 else
"110111011111" when X = 129 AND Y = 125 else
"110111011111" when X = 130 AND Y = 125 else
"110111011111" when X = 131 AND Y = 125 else
"110111011111" when X = 132 AND Y = 125 else
"110111011111" when X = 133 AND Y = 125 else
"110111011111" when X = 134 AND Y = 125 else
"110111011111" when X = 135 AND Y = 125 else
"110111011111" when X = 136 AND Y = 125 else
"110111011111" when X = 137 AND Y = 125 else
"110111011111" when X = 138 AND Y = 125 else
"110111011111" when X = 139 AND Y = 125 else
"110111011111" when X = 140 AND Y = 125 else
"110111011111" when X = 141 AND Y = 125 else
"110111011111" when X = 142 AND Y = 125 else
"110111011111" when X = 143 AND Y = 125 else
"110111011111" when X = 144 AND Y = 125 else
"110111011111" when X = 145 AND Y = 125 else
"110111011111" when X = 146 AND Y = 125 else
"110111011111" when X = 147 AND Y = 125 else
"110111011111" when X = 148 AND Y = 125 else
"110111011111" when X = 149 AND Y = 125 else
"110111011111" when X = 150 AND Y = 125 else
"110111011111" when X = 151 AND Y = 125 else
"110111011111" when X = 152 AND Y = 125 else
"110111011111" when X = 153 AND Y = 125 else
"110111011111" when X = 154 AND Y = 125 else
"110111011111" when X = 155 AND Y = 125 else
"110111011111" when X = 156 AND Y = 125 else
"110111011111" when X = 157 AND Y = 125 else
"110111011111" when X = 158 AND Y = 125 else
"110111011111" when X = 159 AND Y = 125 else
"110111011111" when X = 160 AND Y = 125 else
"110111011111" when X = 161 AND Y = 125 else
"110111011111" when X = 162 AND Y = 125 else
"110111011111" when X = 163 AND Y = 125 else
"110111011111" when X = 164 AND Y = 125 else
"110111011111" when X = 165 AND Y = 125 else
"110111011111" when X = 166 AND Y = 125 else
"110111011111" when X = 167 AND Y = 125 else
"110111011111" when X = 168 AND Y = 125 else
"110111011111" when X = 169 AND Y = 125 else
"110111011111" when X = 170 AND Y = 125 else
"110111011111" when X = 171 AND Y = 125 else
"110111011111" when X = 172 AND Y = 125 else
"110111011111" when X = 173 AND Y = 125 else
"110111011111" when X = 174 AND Y = 125 else
"110111011111" when X = 175 AND Y = 125 else
"110111011111" when X = 176 AND Y = 125 else
"110111011111" when X = 177 AND Y = 125 else
"110111011111" when X = 178 AND Y = 125 else
"110111011111" when X = 179 AND Y = 125 else
"110111011111" when X = 180 AND Y = 125 else
"110111011111" when X = 181 AND Y = 125 else
"110111011111" when X = 182 AND Y = 125 else
"110111011111" when X = 183 AND Y = 125 else
"110111011111" when X = 184 AND Y = 125 else
"110111011111" when X = 185 AND Y = 125 else
"110111011111" when X = 186 AND Y = 125 else
"110111011111" when X = 187 AND Y = 125 else
"110111011111" when X = 188 AND Y = 125 else
"110111011111" when X = 189 AND Y = 125 else
"110111011111" when X = 190 AND Y = 125 else
"110111011111" when X = 191 AND Y = 125 else
"110111011111" when X = 192 AND Y = 125 else
"110111011111" when X = 193 AND Y = 125 else
"110111011111" when X = 194 AND Y = 125 else
"110111011111" when X = 195 AND Y = 125 else
"110111011111" when X = 196 AND Y = 125 else
"110111011111" when X = 197 AND Y = 125 else
"110111011111" when X = 198 AND Y = 125 else
"110111011111" when X = 199 AND Y = 125 else
"110111011111" when X = 200 AND Y = 125 else
"110111011111" when X = 201 AND Y = 125 else
"110111011111" when X = 202 AND Y = 125 else
"110111011111" when X = 203 AND Y = 125 else
"110111011111" when X = 204 AND Y = 125 else
"110111011111" when X = 205 AND Y = 125 else
"110111011111" when X = 206 AND Y = 125 else
"110111011111" when X = 207 AND Y = 125 else
"110111011111" when X = 208 AND Y = 125 else
"110111011111" when X = 209 AND Y = 125 else
"110111011111" when X = 210 AND Y = 125 else
"110111011111" when X = 211 AND Y = 125 else
"110111011111" when X = 212 AND Y = 125 else
"110111011111" when X = 213 AND Y = 125 else
"110111011111" when X = 214 AND Y = 125 else
"110111011111" when X = 215 AND Y = 125 else
"110111011111" when X = 216 AND Y = 125 else
"110111011111" when X = 217 AND Y = 125 else
"110111011111" when X = 218 AND Y = 125 else
"110111011111" when X = 219 AND Y = 125 else
"110111011111" when X = 220 AND Y = 125 else
"110111011111" when X = 221 AND Y = 125 else
"110111011111" when X = 222 AND Y = 125 else
"110111011111" when X = 223 AND Y = 125 else
"110111011111" when X = 224 AND Y = 125 else
"110111011111" when X = 225 AND Y = 125 else
"110111011111" when X = 226 AND Y = 125 else
"110111011111" when X = 227 AND Y = 125 else
"110111011111" when X = 228 AND Y = 125 else
"110111011111" when X = 229 AND Y = 125 else
"110111011111" when X = 230 AND Y = 125 else
"110111011111" when X = 231 AND Y = 125 else
"110111011111" when X = 232 AND Y = 125 else
"110111011111" when X = 233 AND Y = 125 else
"110111011111" when X = 234 AND Y = 125 else
"000000000000" when X = 235 AND Y = 125 else
"000000000000" when X = 236 AND Y = 125 else
"000000000000" when X = 237 AND Y = 125 else
"000000000000" when X = 238 AND Y = 125 else
"000000000000" when X = 239 AND Y = 125 else
"000000000000" when X = 240 AND Y = 125 else
"000000000000" when X = 241 AND Y = 125 else
"000000000000" when X = 242 AND Y = 125 else
"000000000000" when X = 243 AND Y = 125 else
"000000000000" when X = 244 AND Y = 125 else
"110111011111" when X = 245 AND Y = 125 else
"110111011111" when X = 246 AND Y = 125 else
"110111011111" when X = 247 AND Y = 125 else
"110111011111" when X = 248 AND Y = 125 else
"110111011111" when X = 249 AND Y = 125 else
"110111011111" when X = 250 AND Y = 125 else
"110111011111" when X = 251 AND Y = 125 else
"110111011111" when X = 252 AND Y = 125 else
"110111011111" when X = 253 AND Y = 125 else
"110111011111" when X = 254 AND Y = 125 else
"110111011111" when X = 255 AND Y = 125 else
"110111011111" when X = 256 AND Y = 125 else
"110111011111" when X = 257 AND Y = 125 else
"110111011111" when X = 258 AND Y = 125 else
"110111011111" when X = 259 AND Y = 125 else
"110111011111" when X = 260 AND Y = 125 else
"110111011111" when X = 261 AND Y = 125 else
"110111011111" when X = 262 AND Y = 125 else
"110111011111" when X = 263 AND Y = 125 else
"110111011111" when X = 264 AND Y = 125 else
"110111011111" when X = 265 AND Y = 125 else
"110111011111" when X = 266 AND Y = 125 else
"110111011111" when X = 267 AND Y = 125 else
"110111011111" when X = 268 AND Y = 125 else
"110111011111" when X = 269 AND Y = 125 else
"110111011111" when X = 270 AND Y = 125 else
"110111011111" when X = 271 AND Y = 125 else
"110111011111" when X = 272 AND Y = 125 else
"110111011111" when X = 273 AND Y = 125 else
"110111011111" when X = 274 AND Y = 125 else
"110111011111" when X = 275 AND Y = 125 else
"110111011111" when X = 276 AND Y = 125 else
"110111011111" when X = 277 AND Y = 125 else
"110111011111" when X = 278 AND Y = 125 else
"110111011111" when X = 279 AND Y = 125 else
"110111011111" when X = 280 AND Y = 125 else
"110111011111" when X = 281 AND Y = 125 else
"110111011111" when X = 282 AND Y = 125 else
"110111011111" when X = 283 AND Y = 125 else
"110111011111" when X = 284 AND Y = 125 else
"110111011111" when X = 285 AND Y = 125 else
"110111011111" when X = 286 AND Y = 125 else
"110111011111" when X = 287 AND Y = 125 else
"110111011111" when X = 288 AND Y = 125 else
"110111011111" when X = 289 AND Y = 125 else
"110111011111" when X = 290 AND Y = 125 else
"110111011111" when X = 291 AND Y = 125 else
"110111011111" when X = 292 AND Y = 125 else
"110111011111" when X = 293 AND Y = 125 else
"110111011111" when X = 294 AND Y = 125 else
"110111011111" when X = 295 AND Y = 125 else
"110111011111" when X = 296 AND Y = 125 else
"110111011111" when X = 297 AND Y = 125 else
"110111011111" when X = 298 AND Y = 125 else
"110111011111" when X = 299 AND Y = 125 else
"110111011111" when X = 300 AND Y = 125 else
"110111011111" when X = 301 AND Y = 125 else
"110111011111" when X = 302 AND Y = 125 else
"110111011111" when X = 303 AND Y = 125 else
"110111011111" when X = 304 AND Y = 125 else
"110111011111" when X = 305 AND Y = 125 else
"110111011111" when X = 306 AND Y = 125 else
"110111011111" when X = 307 AND Y = 125 else
"110111011111" when X = 308 AND Y = 125 else
"110111011111" when X = 309 AND Y = 125 else
"110111011111" when X = 310 AND Y = 125 else
"110111011111" when X = 311 AND Y = 125 else
"110111011111" when X = 312 AND Y = 125 else
"110111011111" when X = 313 AND Y = 125 else
"110111011111" when X = 314 AND Y = 125 else
"110111011111" when X = 315 AND Y = 125 else
"110111011111" when X = 316 AND Y = 125 else
"110111011111" when X = 317 AND Y = 125 else
"110111011111" when X = 318 AND Y = 125 else
"110111011111" when X = 319 AND Y = 125 else
"000000000000" when X = 320 AND Y = 125 else
"000000000000" when X = 321 AND Y = 125 else
"000000000000" when X = 322 AND Y = 125 else
"000000000000" when X = 323 AND Y = 125 else
"000000000000" when X = 324 AND Y = 125 else
"100010011101" when X = 0 AND Y = 126 else
"100010011101" when X = 1 AND Y = 126 else
"100010011101" when X = 2 AND Y = 126 else
"100010011101" when X = 3 AND Y = 126 else
"100010011101" when X = 4 AND Y = 126 else
"100010011101" when X = 5 AND Y = 126 else
"100010011101" when X = 6 AND Y = 126 else
"100010011101" when X = 7 AND Y = 126 else
"100010011101" when X = 8 AND Y = 126 else
"100010011101" when X = 9 AND Y = 126 else
"100010011101" when X = 10 AND Y = 126 else
"100010011101" when X = 11 AND Y = 126 else
"100010011101" when X = 12 AND Y = 126 else
"100010011101" when X = 13 AND Y = 126 else
"100010011101" when X = 14 AND Y = 126 else
"100010011101" when X = 15 AND Y = 126 else
"100010011101" when X = 16 AND Y = 126 else
"100010011101" when X = 17 AND Y = 126 else
"100010011101" when X = 18 AND Y = 126 else
"100010011101" when X = 19 AND Y = 126 else
"100010011101" when X = 20 AND Y = 126 else
"100010011101" when X = 21 AND Y = 126 else
"100010011101" when X = 22 AND Y = 126 else
"100010011101" when X = 23 AND Y = 126 else
"100010011101" when X = 24 AND Y = 126 else
"100010011101" when X = 25 AND Y = 126 else
"100010011101" when X = 26 AND Y = 126 else
"100010011101" when X = 27 AND Y = 126 else
"100010011101" when X = 28 AND Y = 126 else
"100010011101" when X = 29 AND Y = 126 else
"100010011101" when X = 30 AND Y = 126 else
"100010011101" when X = 31 AND Y = 126 else
"100010011101" when X = 32 AND Y = 126 else
"100010011101" when X = 33 AND Y = 126 else
"100010011101" when X = 34 AND Y = 126 else
"100010011101" when X = 35 AND Y = 126 else
"100010011101" when X = 36 AND Y = 126 else
"100010011101" when X = 37 AND Y = 126 else
"100010011101" when X = 38 AND Y = 126 else
"100010011101" when X = 39 AND Y = 126 else
"100010011101" when X = 40 AND Y = 126 else
"100010011101" when X = 41 AND Y = 126 else
"100010011101" when X = 42 AND Y = 126 else
"100010011101" when X = 43 AND Y = 126 else
"100010011101" when X = 44 AND Y = 126 else
"100010011101" when X = 45 AND Y = 126 else
"100010011101" when X = 46 AND Y = 126 else
"100010011101" when X = 47 AND Y = 126 else
"100010011101" when X = 48 AND Y = 126 else
"100010011101" when X = 49 AND Y = 126 else
"100010011101" when X = 50 AND Y = 126 else
"100010011101" when X = 51 AND Y = 126 else
"100010011101" when X = 52 AND Y = 126 else
"100010011101" when X = 53 AND Y = 126 else
"100010011101" when X = 54 AND Y = 126 else
"100010011101" when X = 55 AND Y = 126 else
"100010011101" when X = 56 AND Y = 126 else
"100010011101" when X = 57 AND Y = 126 else
"100010011101" when X = 58 AND Y = 126 else
"100010011101" when X = 59 AND Y = 126 else
"100010011101" when X = 60 AND Y = 126 else
"100010011101" when X = 61 AND Y = 126 else
"100010011101" when X = 62 AND Y = 126 else
"100010011101" when X = 63 AND Y = 126 else
"100010011101" when X = 64 AND Y = 126 else
"100010011101" when X = 65 AND Y = 126 else
"100010011101" when X = 66 AND Y = 126 else
"100010011101" when X = 67 AND Y = 126 else
"100010011101" when X = 68 AND Y = 126 else
"100010011101" when X = 69 AND Y = 126 else
"100010011101" when X = 70 AND Y = 126 else
"100010011101" when X = 71 AND Y = 126 else
"100010011101" when X = 72 AND Y = 126 else
"100010011101" when X = 73 AND Y = 126 else
"100010011101" when X = 74 AND Y = 126 else
"100010011101" when X = 75 AND Y = 126 else
"100010011101" when X = 76 AND Y = 126 else
"100010011101" when X = 77 AND Y = 126 else
"100010011101" when X = 78 AND Y = 126 else
"100010011101" when X = 79 AND Y = 126 else
"100010011101" when X = 80 AND Y = 126 else
"100010011101" when X = 81 AND Y = 126 else
"100010011101" when X = 82 AND Y = 126 else
"100010011101" when X = 83 AND Y = 126 else
"100010011101" when X = 84 AND Y = 126 else
"100010011101" when X = 85 AND Y = 126 else
"100010011101" when X = 86 AND Y = 126 else
"100010011101" when X = 87 AND Y = 126 else
"100010011101" when X = 88 AND Y = 126 else
"100010011101" when X = 89 AND Y = 126 else
"100010011101" when X = 90 AND Y = 126 else
"100010011101" when X = 91 AND Y = 126 else
"100010011101" when X = 92 AND Y = 126 else
"100010011101" when X = 93 AND Y = 126 else
"100010011101" when X = 94 AND Y = 126 else
"100010011101" when X = 95 AND Y = 126 else
"100010011101" when X = 96 AND Y = 126 else
"100010011101" when X = 97 AND Y = 126 else
"100010011101" when X = 98 AND Y = 126 else
"100010011101" when X = 99 AND Y = 126 else
"100010011101" when X = 100 AND Y = 126 else
"100010011101" when X = 101 AND Y = 126 else
"100010011101" when X = 102 AND Y = 126 else
"100010011101" when X = 103 AND Y = 126 else
"100010011101" when X = 104 AND Y = 126 else
"100010011101" when X = 105 AND Y = 126 else
"100010011101" when X = 106 AND Y = 126 else
"100010011101" when X = 107 AND Y = 126 else
"100010011101" when X = 108 AND Y = 126 else
"100010011101" when X = 109 AND Y = 126 else
"110111011111" when X = 110 AND Y = 126 else
"110111011111" when X = 111 AND Y = 126 else
"110111011111" when X = 112 AND Y = 126 else
"110111011111" when X = 113 AND Y = 126 else
"110111011111" when X = 114 AND Y = 126 else
"110111011111" when X = 115 AND Y = 126 else
"110111011111" when X = 116 AND Y = 126 else
"110111011111" when X = 117 AND Y = 126 else
"110111011111" when X = 118 AND Y = 126 else
"110111011111" when X = 119 AND Y = 126 else
"110111011111" when X = 120 AND Y = 126 else
"110111011111" when X = 121 AND Y = 126 else
"110111011111" when X = 122 AND Y = 126 else
"110111011111" when X = 123 AND Y = 126 else
"110111011111" when X = 124 AND Y = 126 else
"110111011111" when X = 125 AND Y = 126 else
"110111011111" when X = 126 AND Y = 126 else
"110111011111" when X = 127 AND Y = 126 else
"110111011111" when X = 128 AND Y = 126 else
"110111011111" when X = 129 AND Y = 126 else
"110111011111" when X = 130 AND Y = 126 else
"110111011111" when X = 131 AND Y = 126 else
"110111011111" when X = 132 AND Y = 126 else
"110111011111" when X = 133 AND Y = 126 else
"110111011111" when X = 134 AND Y = 126 else
"110111011111" when X = 135 AND Y = 126 else
"110111011111" when X = 136 AND Y = 126 else
"110111011111" when X = 137 AND Y = 126 else
"110111011111" when X = 138 AND Y = 126 else
"110111011111" when X = 139 AND Y = 126 else
"110111011111" when X = 140 AND Y = 126 else
"110111011111" when X = 141 AND Y = 126 else
"110111011111" when X = 142 AND Y = 126 else
"110111011111" when X = 143 AND Y = 126 else
"110111011111" when X = 144 AND Y = 126 else
"110111011111" when X = 145 AND Y = 126 else
"110111011111" when X = 146 AND Y = 126 else
"110111011111" when X = 147 AND Y = 126 else
"110111011111" when X = 148 AND Y = 126 else
"110111011111" when X = 149 AND Y = 126 else
"110111011111" when X = 150 AND Y = 126 else
"110111011111" when X = 151 AND Y = 126 else
"110111011111" when X = 152 AND Y = 126 else
"110111011111" when X = 153 AND Y = 126 else
"110111011111" when X = 154 AND Y = 126 else
"110111011111" when X = 155 AND Y = 126 else
"110111011111" when X = 156 AND Y = 126 else
"110111011111" when X = 157 AND Y = 126 else
"110111011111" when X = 158 AND Y = 126 else
"110111011111" when X = 159 AND Y = 126 else
"110111011111" when X = 160 AND Y = 126 else
"110111011111" when X = 161 AND Y = 126 else
"110111011111" when X = 162 AND Y = 126 else
"110111011111" when X = 163 AND Y = 126 else
"110111011111" when X = 164 AND Y = 126 else
"110111011111" when X = 165 AND Y = 126 else
"110111011111" when X = 166 AND Y = 126 else
"110111011111" when X = 167 AND Y = 126 else
"110111011111" when X = 168 AND Y = 126 else
"110111011111" when X = 169 AND Y = 126 else
"110111011111" when X = 170 AND Y = 126 else
"110111011111" when X = 171 AND Y = 126 else
"110111011111" when X = 172 AND Y = 126 else
"110111011111" when X = 173 AND Y = 126 else
"110111011111" when X = 174 AND Y = 126 else
"110111011111" when X = 175 AND Y = 126 else
"110111011111" when X = 176 AND Y = 126 else
"110111011111" when X = 177 AND Y = 126 else
"110111011111" when X = 178 AND Y = 126 else
"110111011111" when X = 179 AND Y = 126 else
"110111011111" when X = 180 AND Y = 126 else
"110111011111" when X = 181 AND Y = 126 else
"110111011111" when X = 182 AND Y = 126 else
"110111011111" when X = 183 AND Y = 126 else
"110111011111" when X = 184 AND Y = 126 else
"110111011111" when X = 185 AND Y = 126 else
"110111011111" when X = 186 AND Y = 126 else
"110111011111" when X = 187 AND Y = 126 else
"110111011111" when X = 188 AND Y = 126 else
"110111011111" when X = 189 AND Y = 126 else
"110111011111" when X = 190 AND Y = 126 else
"110111011111" when X = 191 AND Y = 126 else
"110111011111" when X = 192 AND Y = 126 else
"110111011111" when X = 193 AND Y = 126 else
"110111011111" when X = 194 AND Y = 126 else
"110111011111" when X = 195 AND Y = 126 else
"110111011111" when X = 196 AND Y = 126 else
"110111011111" when X = 197 AND Y = 126 else
"110111011111" when X = 198 AND Y = 126 else
"110111011111" when X = 199 AND Y = 126 else
"110111011111" when X = 200 AND Y = 126 else
"110111011111" when X = 201 AND Y = 126 else
"110111011111" when X = 202 AND Y = 126 else
"110111011111" when X = 203 AND Y = 126 else
"110111011111" when X = 204 AND Y = 126 else
"110111011111" when X = 205 AND Y = 126 else
"110111011111" when X = 206 AND Y = 126 else
"110111011111" when X = 207 AND Y = 126 else
"110111011111" when X = 208 AND Y = 126 else
"110111011111" when X = 209 AND Y = 126 else
"110111011111" when X = 210 AND Y = 126 else
"110111011111" when X = 211 AND Y = 126 else
"110111011111" when X = 212 AND Y = 126 else
"110111011111" when X = 213 AND Y = 126 else
"110111011111" when X = 214 AND Y = 126 else
"110111011111" when X = 215 AND Y = 126 else
"110111011111" when X = 216 AND Y = 126 else
"110111011111" when X = 217 AND Y = 126 else
"110111011111" when X = 218 AND Y = 126 else
"110111011111" when X = 219 AND Y = 126 else
"110111011111" when X = 220 AND Y = 126 else
"110111011111" when X = 221 AND Y = 126 else
"110111011111" when X = 222 AND Y = 126 else
"110111011111" when X = 223 AND Y = 126 else
"110111011111" when X = 224 AND Y = 126 else
"110111011111" when X = 225 AND Y = 126 else
"110111011111" when X = 226 AND Y = 126 else
"110111011111" when X = 227 AND Y = 126 else
"110111011111" when X = 228 AND Y = 126 else
"110111011111" when X = 229 AND Y = 126 else
"110111011111" when X = 230 AND Y = 126 else
"110111011111" when X = 231 AND Y = 126 else
"110111011111" when X = 232 AND Y = 126 else
"110111011111" when X = 233 AND Y = 126 else
"110111011111" when X = 234 AND Y = 126 else
"000000000000" when X = 235 AND Y = 126 else
"000000000000" when X = 236 AND Y = 126 else
"000000000000" when X = 237 AND Y = 126 else
"000000000000" when X = 238 AND Y = 126 else
"000000000000" when X = 239 AND Y = 126 else
"000000000000" when X = 240 AND Y = 126 else
"000000000000" when X = 241 AND Y = 126 else
"000000000000" when X = 242 AND Y = 126 else
"000000000000" when X = 243 AND Y = 126 else
"000000000000" when X = 244 AND Y = 126 else
"110111011111" when X = 245 AND Y = 126 else
"110111011111" when X = 246 AND Y = 126 else
"110111011111" when X = 247 AND Y = 126 else
"110111011111" when X = 248 AND Y = 126 else
"110111011111" when X = 249 AND Y = 126 else
"110111011111" when X = 250 AND Y = 126 else
"110111011111" when X = 251 AND Y = 126 else
"110111011111" when X = 252 AND Y = 126 else
"110111011111" when X = 253 AND Y = 126 else
"110111011111" when X = 254 AND Y = 126 else
"110111011111" when X = 255 AND Y = 126 else
"110111011111" when X = 256 AND Y = 126 else
"110111011111" when X = 257 AND Y = 126 else
"110111011111" when X = 258 AND Y = 126 else
"110111011111" when X = 259 AND Y = 126 else
"110111011111" when X = 260 AND Y = 126 else
"110111011111" when X = 261 AND Y = 126 else
"110111011111" when X = 262 AND Y = 126 else
"110111011111" when X = 263 AND Y = 126 else
"110111011111" when X = 264 AND Y = 126 else
"110111011111" when X = 265 AND Y = 126 else
"110111011111" when X = 266 AND Y = 126 else
"110111011111" when X = 267 AND Y = 126 else
"110111011111" when X = 268 AND Y = 126 else
"110111011111" when X = 269 AND Y = 126 else
"110111011111" when X = 270 AND Y = 126 else
"110111011111" when X = 271 AND Y = 126 else
"110111011111" when X = 272 AND Y = 126 else
"110111011111" when X = 273 AND Y = 126 else
"110111011111" when X = 274 AND Y = 126 else
"110111011111" when X = 275 AND Y = 126 else
"110111011111" when X = 276 AND Y = 126 else
"110111011111" when X = 277 AND Y = 126 else
"110111011111" when X = 278 AND Y = 126 else
"110111011111" when X = 279 AND Y = 126 else
"110111011111" when X = 280 AND Y = 126 else
"110111011111" when X = 281 AND Y = 126 else
"110111011111" when X = 282 AND Y = 126 else
"110111011111" when X = 283 AND Y = 126 else
"110111011111" when X = 284 AND Y = 126 else
"110111011111" when X = 285 AND Y = 126 else
"110111011111" when X = 286 AND Y = 126 else
"110111011111" when X = 287 AND Y = 126 else
"110111011111" when X = 288 AND Y = 126 else
"110111011111" when X = 289 AND Y = 126 else
"110111011111" when X = 290 AND Y = 126 else
"110111011111" when X = 291 AND Y = 126 else
"110111011111" when X = 292 AND Y = 126 else
"110111011111" when X = 293 AND Y = 126 else
"110111011111" when X = 294 AND Y = 126 else
"110111011111" when X = 295 AND Y = 126 else
"110111011111" when X = 296 AND Y = 126 else
"110111011111" when X = 297 AND Y = 126 else
"110111011111" when X = 298 AND Y = 126 else
"110111011111" when X = 299 AND Y = 126 else
"110111011111" when X = 300 AND Y = 126 else
"110111011111" when X = 301 AND Y = 126 else
"110111011111" when X = 302 AND Y = 126 else
"110111011111" when X = 303 AND Y = 126 else
"110111011111" when X = 304 AND Y = 126 else
"110111011111" when X = 305 AND Y = 126 else
"110111011111" when X = 306 AND Y = 126 else
"110111011111" when X = 307 AND Y = 126 else
"110111011111" when X = 308 AND Y = 126 else
"110111011111" when X = 309 AND Y = 126 else
"110111011111" when X = 310 AND Y = 126 else
"110111011111" when X = 311 AND Y = 126 else
"110111011111" when X = 312 AND Y = 126 else
"110111011111" when X = 313 AND Y = 126 else
"110111011111" when X = 314 AND Y = 126 else
"110111011111" when X = 315 AND Y = 126 else
"110111011111" when X = 316 AND Y = 126 else
"110111011111" when X = 317 AND Y = 126 else
"110111011111" when X = 318 AND Y = 126 else
"110111011111" when X = 319 AND Y = 126 else
"000000000000" when X = 320 AND Y = 126 else
"000000000000" when X = 321 AND Y = 126 else
"000000000000" when X = 322 AND Y = 126 else
"000000000000" when X = 323 AND Y = 126 else
"000000000000" when X = 324 AND Y = 126 else
"100010011101" when X = 0 AND Y = 127 else
"100010011101" when X = 1 AND Y = 127 else
"100010011101" when X = 2 AND Y = 127 else
"100010011101" when X = 3 AND Y = 127 else
"100010011101" when X = 4 AND Y = 127 else
"100010011101" when X = 5 AND Y = 127 else
"100010011101" when X = 6 AND Y = 127 else
"100010011101" when X = 7 AND Y = 127 else
"100010011101" when X = 8 AND Y = 127 else
"100010011101" when X = 9 AND Y = 127 else
"100010011101" when X = 10 AND Y = 127 else
"100010011101" when X = 11 AND Y = 127 else
"100010011101" when X = 12 AND Y = 127 else
"100010011101" when X = 13 AND Y = 127 else
"100010011101" when X = 14 AND Y = 127 else
"100010011101" when X = 15 AND Y = 127 else
"100010011101" when X = 16 AND Y = 127 else
"100010011101" when X = 17 AND Y = 127 else
"100010011101" when X = 18 AND Y = 127 else
"100010011101" when X = 19 AND Y = 127 else
"100010011101" when X = 20 AND Y = 127 else
"100010011101" when X = 21 AND Y = 127 else
"100010011101" when X = 22 AND Y = 127 else
"100010011101" when X = 23 AND Y = 127 else
"100010011101" when X = 24 AND Y = 127 else
"100010011101" when X = 25 AND Y = 127 else
"100010011101" when X = 26 AND Y = 127 else
"100010011101" when X = 27 AND Y = 127 else
"100010011101" when X = 28 AND Y = 127 else
"100010011101" when X = 29 AND Y = 127 else
"100010011101" when X = 30 AND Y = 127 else
"100010011101" when X = 31 AND Y = 127 else
"100010011101" when X = 32 AND Y = 127 else
"100010011101" when X = 33 AND Y = 127 else
"100010011101" when X = 34 AND Y = 127 else
"100010011101" when X = 35 AND Y = 127 else
"100010011101" when X = 36 AND Y = 127 else
"100010011101" when X = 37 AND Y = 127 else
"100010011101" when X = 38 AND Y = 127 else
"100010011101" when X = 39 AND Y = 127 else
"100010011101" when X = 40 AND Y = 127 else
"100010011101" when X = 41 AND Y = 127 else
"100010011101" when X = 42 AND Y = 127 else
"100010011101" when X = 43 AND Y = 127 else
"100010011101" when X = 44 AND Y = 127 else
"100010011101" when X = 45 AND Y = 127 else
"100010011101" when X = 46 AND Y = 127 else
"100010011101" when X = 47 AND Y = 127 else
"100010011101" when X = 48 AND Y = 127 else
"100010011101" when X = 49 AND Y = 127 else
"100010011101" when X = 50 AND Y = 127 else
"100010011101" when X = 51 AND Y = 127 else
"100010011101" when X = 52 AND Y = 127 else
"100010011101" when X = 53 AND Y = 127 else
"100010011101" when X = 54 AND Y = 127 else
"100010011101" when X = 55 AND Y = 127 else
"100010011101" when X = 56 AND Y = 127 else
"100010011101" when X = 57 AND Y = 127 else
"100010011101" when X = 58 AND Y = 127 else
"100010011101" when X = 59 AND Y = 127 else
"100010011101" when X = 60 AND Y = 127 else
"100010011101" when X = 61 AND Y = 127 else
"100010011101" when X = 62 AND Y = 127 else
"100010011101" when X = 63 AND Y = 127 else
"100010011101" when X = 64 AND Y = 127 else
"100010011101" when X = 65 AND Y = 127 else
"100010011101" when X = 66 AND Y = 127 else
"100010011101" when X = 67 AND Y = 127 else
"100010011101" when X = 68 AND Y = 127 else
"100010011101" when X = 69 AND Y = 127 else
"100010011101" when X = 70 AND Y = 127 else
"100010011101" when X = 71 AND Y = 127 else
"100010011101" when X = 72 AND Y = 127 else
"100010011101" when X = 73 AND Y = 127 else
"100010011101" when X = 74 AND Y = 127 else
"100010011101" when X = 75 AND Y = 127 else
"100010011101" when X = 76 AND Y = 127 else
"100010011101" when X = 77 AND Y = 127 else
"100010011101" when X = 78 AND Y = 127 else
"100010011101" when X = 79 AND Y = 127 else
"100010011101" when X = 80 AND Y = 127 else
"100010011101" when X = 81 AND Y = 127 else
"100010011101" when X = 82 AND Y = 127 else
"100010011101" when X = 83 AND Y = 127 else
"100010011101" when X = 84 AND Y = 127 else
"100010011101" when X = 85 AND Y = 127 else
"100010011101" when X = 86 AND Y = 127 else
"100010011101" when X = 87 AND Y = 127 else
"100010011101" when X = 88 AND Y = 127 else
"100010011101" when X = 89 AND Y = 127 else
"100010011101" when X = 90 AND Y = 127 else
"100010011101" when X = 91 AND Y = 127 else
"100010011101" when X = 92 AND Y = 127 else
"100010011101" when X = 93 AND Y = 127 else
"100010011101" when X = 94 AND Y = 127 else
"100010011101" when X = 95 AND Y = 127 else
"100010011101" when X = 96 AND Y = 127 else
"100010011101" when X = 97 AND Y = 127 else
"100010011101" when X = 98 AND Y = 127 else
"100010011101" when X = 99 AND Y = 127 else
"100010011101" when X = 100 AND Y = 127 else
"100010011101" when X = 101 AND Y = 127 else
"100010011101" when X = 102 AND Y = 127 else
"100010011101" when X = 103 AND Y = 127 else
"100010011101" when X = 104 AND Y = 127 else
"100010011101" when X = 105 AND Y = 127 else
"100010011101" when X = 106 AND Y = 127 else
"100010011101" when X = 107 AND Y = 127 else
"100010011101" when X = 108 AND Y = 127 else
"100010011101" when X = 109 AND Y = 127 else
"110111011111" when X = 110 AND Y = 127 else
"110111011111" when X = 111 AND Y = 127 else
"110111011111" when X = 112 AND Y = 127 else
"110111011111" when X = 113 AND Y = 127 else
"110111011111" when X = 114 AND Y = 127 else
"110111011111" when X = 115 AND Y = 127 else
"110111011111" when X = 116 AND Y = 127 else
"110111011111" when X = 117 AND Y = 127 else
"110111011111" when X = 118 AND Y = 127 else
"110111011111" when X = 119 AND Y = 127 else
"110111011111" when X = 120 AND Y = 127 else
"110111011111" when X = 121 AND Y = 127 else
"110111011111" when X = 122 AND Y = 127 else
"110111011111" when X = 123 AND Y = 127 else
"110111011111" when X = 124 AND Y = 127 else
"110111011111" when X = 125 AND Y = 127 else
"110111011111" when X = 126 AND Y = 127 else
"110111011111" when X = 127 AND Y = 127 else
"110111011111" when X = 128 AND Y = 127 else
"110111011111" when X = 129 AND Y = 127 else
"110111011111" when X = 130 AND Y = 127 else
"110111011111" when X = 131 AND Y = 127 else
"110111011111" when X = 132 AND Y = 127 else
"110111011111" when X = 133 AND Y = 127 else
"110111011111" when X = 134 AND Y = 127 else
"110111011111" when X = 135 AND Y = 127 else
"110111011111" when X = 136 AND Y = 127 else
"110111011111" when X = 137 AND Y = 127 else
"110111011111" when X = 138 AND Y = 127 else
"110111011111" when X = 139 AND Y = 127 else
"110111011111" when X = 140 AND Y = 127 else
"110111011111" when X = 141 AND Y = 127 else
"110111011111" when X = 142 AND Y = 127 else
"110111011111" when X = 143 AND Y = 127 else
"110111011111" when X = 144 AND Y = 127 else
"110111011111" when X = 145 AND Y = 127 else
"110111011111" when X = 146 AND Y = 127 else
"110111011111" when X = 147 AND Y = 127 else
"110111011111" when X = 148 AND Y = 127 else
"110111011111" when X = 149 AND Y = 127 else
"110111011111" when X = 150 AND Y = 127 else
"110111011111" when X = 151 AND Y = 127 else
"110111011111" when X = 152 AND Y = 127 else
"110111011111" when X = 153 AND Y = 127 else
"110111011111" when X = 154 AND Y = 127 else
"110111011111" when X = 155 AND Y = 127 else
"110111011111" when X = 156 AND Y = 127 else
"110111011111" when X = 157 AND Y = 127 else
"110111011111" when X = 158 AND Y = 127 else
"110111011111" when X = 159 AND Y = 127 else
"110111011111" when X = 160 AND Y = 127 else
"110111011111" when X = 161 AND Y = 127 else
"110111011111" when X = 162 AND Y = 127 else
"110111011111" when X = 163 AND Y = 127 else
"110111011111" when X = 164 AND Y = 127 else
"110111011111" when X = 165 AND Y = 127 else
"110111011111" when X = 166 AND Y = 127 else
"110111011111" when X = 167 AND Y = 127 else
"110111011111" when X = 168 AND Y = 127 else
"110111011111" when X = 169 AND Y = 127 else
"110111011111" when X = 170 AND Y = 127 else
"110111011111" when X = 171 AND Y = 127 else
"110111011111" when X = 172 AND Y = 127 else
"110111011111" when X = 173 AND Y = 127 else
"110111011111" when X = 174 AND Y = 127 else
"110111011111" when X = 175 AND Y = 127 else
"110111011111" when X = 176 AND Y = 127 else
"110111011111" when X = 177 AND Y = 127 else
"110111011111" when X = 178 AND Y = 127 else
"110111011111" when X = 179 AND Y = 127 else
"110111011111" when X = 180 AND Y = 127 else
"110111011111" when X = 181 AND Y = 127 else
"110111011111" when X = 182 AND Y = 127 else
"110111011111" when X = 183 AND Y = 127 else
"110111011111" when X = 184 AND Y = 127 else
"110111011111" when X = 185 AND Y = 127 else
"110111011111" when X = 186 AND Y = 127 else
"110111011111" when X = 187 AND Y = 127 else
"110111011111" when X = 188 AND Y = 127 else
"110111011111" when X = 189 AND Y = 127 else
"110111011111" when X = 190 AND Y = 127 else
"110111011111" when X = 191 AND Y = 127 else
"110111011111" when X = 192 AND Y = 127 else
"110111011111" when X = 193 AND Y = 127 else
"110111011111" when X = 194 AND Y = 127 else
"110111011111" when X = 195 AND Y = 127 else
"110111011111" when X = 196 AND Y = 127 else
"110111011111" when X = 197 AND Y = 127 else
"110111011111" when X = 198 AND Y = 127 else
"110111011111" when X = 199 AND Y = 127 else
"110111011111" when X = 200 AND Y = 127 else
"110111011111" when X = 201 AND Y = 127 else
"110111011111" when X = 202 AND Y = 127 else
"110111011111" when X = 203 AND Y = 127 else
"110111011111" when X = 204 AND Y = 127 else
"110111011111" when X = 205 AND Y = 127 else
"110111011111" when X = 206 AND Y = 127 else
"110111011111" when X = 207 AND Y = 127 else
"110111011111" when X = 208 AND Y = 127 else
"110111011111" when X = 209 AND Y = 127 else
"110111011111" when X = 210 AND Y = 127 else
"110111011111" when X = 211 AND Y = 127 else
"110111011111" when X = 212 AND Y = 127 else
"110111011111" when X = 213 AND Y = 127 else
"110111011111" when X = 214 AND Y = 127 else
"110111011111" when X = 215 AND Y = 127 else
"110111011111" when X = 216 AND Y = 127 else
"110111011111" when X = 217 AND Y = 127 else
"110111011111" when X = 218 AND Y = 127 else
"110111011111" when X = 219 AND Y = 127 else
"110111011111" when X = 220 AND Y = 127 else
"110111011111" when X = 221 AND Y = 127 else
"110111011111" when X = 222 AND Y = 127 else
"110111011111" when X = 223 AND Y = 127 else
"110111011111" when X = 224 AND Y = 127 else
"110111011111" when X = 225 AND Y = 127 else
"110111011111" when X = 226 AND Y = 127 else
"110111011111" when X = 227 AND Y = 127 else
"110111011111" when X = 228 AND Y = 127 else
"110111011111" when X = 229 AND Y = 127 else
"110111011111" when X = 230 AND Y = 127 else
"110111011111" when X = 231 AND Y = 127 else
"110111011111" when X = 232 AND Y = 127 else
"110111011111" when X = 233 AND Y = 127 else
"110111011111" when X = 234 AND Y = 127 else
"000000000000" when X = 235 AND Y = 127 else
"000000000000" when X = 236 AND Y = 127 else
"000000000000" when X = 237 AND Y = 127 else
"000000000000" when X = 238 AND Y = 127 else
"000000000000" when X = 239 AND Y = 127 else
"000000000000" when X = 240 AND Y = 127 else
"000000000000" when X = 241 AND Y = 127 else
"000000000000" when X = 242 AND Y = 127 else
"000000000000" when X = 243 AND Y = 127 else
"000000000000" when X = 244 AND Y = 127 else
"110111011111" when X = 245 AND Y = 127 else
"110111011111" when X = 246 AND Y = 127 else
"110111011111" when X = 247 AND Y = 127 else
"110111011111" when X = 248 AND Y = 127 else
"110111011111" when X = 249 AND Y = 127 else
"110111011111" when X = 250 AND Y = 127 else
"110111011111" when X = 251 AND Y = 127 else
"110111011111" when X = 252 AND Y = 127 else
"110111011111" when X = 253 AND Y = 127 else
"110111011111" when X = 254 AND Y = 127 else
"110111011111" when X = 255 AND Y = 127 else
"110111011111" when X = 256 AND Y = 127 else
"110111011111" when X = 257 AND Y = 127 else
"110111011111" when X = 258 AND Y = 127 else
"110111011111" when X = 259 AND Y = 127 else
"110111011111" when X = 260 AND Y = 127 else
"110111011111" when X = 261 AND Y = 127 else
"110111011111" when X = 262 AND Y = 127 else
"110111011111" when X = 263 AND Y = 127 else
"110111011111" when X = 264 AND Y = 127 else
"110111011111" when X = 265 AND Y = 127 else
"110111011111" when X = 266 AND Y = 127 else
"110111011111" when X = 267 AND Y = 127 else
"110111011111" when X = 268 AND Y = 127 else
"110111011111" when X = 269 AND Y = 127 else
"110111011111" when X = 270 AND Y = 127 else
"110111011111" when X = 271 AND Y = 127 else
"110111011111" when X = 272 AND Y = 127 else
"110111011111" when X = 273 AND Y = 127 else
"110111011111" when X = 274 AND Y = 127 else
"110111011111" when X = 275 AND Y = 127 else
"110111011111" when X = 276 AND Y = 127 else
"110111011111" when X = 277 AND Y = 127 else
"110111011111" when X = 278 AND Y = 127 else
"110111011111" when X = 279 AND Y = 127 else
"110111011111" when X = 280 AND Y = 127 else
"110111011111" when X = 281 AND Y = 127 else
"110111011111" when X = 282 AND Y = 127 else
"110111011111" when X = 283 AND Y = 127 else
"110111011111" when X = 284 AND Y = 127 else
"110111011111" when X = 285 AND Y = 127 else
"110111011111" when X = 286 AND Y = 127 else
"110111011111" when X = 287 AND Y = 127 else
"110111011111" when X = 288 AND Y = 127 else
"110111011111" when X = 289 AND Y = 127 else
"110111011111" when X = 290 AND Y = 127 else
"110111011111" when X = 291 AND Y = 127 else
"110111011111" when X = 292 AND Y = 127 else
"110111011111" when X = 293 AND Y = 127 else
"110111011111" when X = 294 AND Y = 127 else
"110111011111" when X = 295 AND Y = 127 else
"110111011111" when X = 296 AND Y = 127 else
"110111011111" when X = 297 AND Y = 127 else
"110111011111" when X = 298 AND Y = 127 else
"110111011111" when X = 299 AND Y = 127 else
"110111011111" when X = 300 AND Y = 127 else
"110111011111" when X = 301 AND Y = 127 else
"110111011111" when X = 302 AND Y = 127 else
"110111011111" when X = 303 AND Y = 127 else
"110111011111" when X = 304 AND Y = 127 else
"110111011111" when X = 305 AND Y = 127 else
"110111011111" when X = 306 AND Y = 127 else
"110111011111" when X = 307 AND Y = 127 else
"110111011111" when X = 308 AND Y = 127 else
"110111011111" when X = 309 AND Y = 127 else
"110111011111" when X = 310 AND Y = 127 else
"110111011111" when X = 311 AND Y = 127 else
"110111011111" when X = 312 AND Y = 127 else
"110111011111" when X = 313 AND Y = 127 else
"110111011111" when X = 314 AND Y = 127 else
"110111011111" when X = 315 AND Y = 127 else
"110111011111" when X = 316 AND Y = 127 else
"110111011111" when X = 317 AND Y = 127 else
"110111011111" when X = 318 AND Y = 127 else
"110111011111" when X = 319 AND Y = 127 else
"000000000000" when X = 320 AND Y = 127 else
"000000000000" when X = 321 AND Y = 127 else
"000000000000" when X = 322 AND Y = 127 else
"000000000000" when X = 323 AND Y = 127 else
"000000000000" when X = 324 AND Y = 127 else
"100010011101" when X = 0 AND Y = 128 else
"100010011101" when X = 1 AND Y = 128 else
"100010011101" when X = 2 AND Y = 128 else
"100010011101" when X = 3 AND Y = 128 else
"100010011101" when X = 4 AND Y = 128 else
"100010011101" when X = 5 AND Y = 128 else
"100010011101" when X = 6 AND Y = 128 else
"100010011101" when X = 7 AND Y = 128 else
"100010011101" when X = 8 AND Y = 128 else
"100010011101" when X = 9 AND Y = 128 else
"100010011101" when X = 10 AND Y = 128 else
"100010011101" when X = 11 AND Y = 128 else
"100010011101" when X = 12 AND Y = 128 else
"100010011101" when X = 13 AND Y = 128 else
"100010011101" when X = 14 AND Y = 128 else
"100010011101" when X = 15 AND Y = 128 else
"100010011101" when X = 16 AND Y = 128 else
"100010011101" when X = 17 AND Y = 128 else
"100010011101" when X = 18 AND Y = 128 else
"100010011101" when X = 19 AND Y = 128 else
"100010011101" when X = 20 AND Y = 128 else
"100010011101" when X = 21 AND Y = 128 else
"100010011101" when X = 22 AND Y = 128 else
"100010011101" when X = 23 AND Y = 128 else
"100010011101" when X = 24 AND Y = 128 else
"100010011101" when X = 25 AND Y = 128 else
"100010011101" when X = 26 AND Y = 128 else
"100010011101" when X = 27 AND Y = 128 else
"100010011101" when X = 28 AND Y = 128 else
"100010011101" when X = 29 AND Y = 128 else
"100010011101" when X = 30 AND Y = 128 else
"100010011101" when X = 31 AND Y = 128 else
"100010011101" when X = 32 AND Y = 128 else
"100010011101" when X = 33 AND Y = 128 else
"100010011101" when X = 34 AND Y = 128 else
"100010011101" when X = 35 AND Y = 128 else
"100010011101" when X = 36 AND Y = 128 else
"100010011101" when X = 37 AND Y = 128 else
"100010011101" when X = 38 AND Y = 128 else
"100010011101" when X = 39 AND Y = 128 else
"100010011101" when X = 40 AND Y = 128 else
"100010011101" when X = 41 AND Y = 128 else
"100010011101" when X = 42 AND Y = 128 else
"100010011101" when X = 43 AND Y = 128 else
"100010011101" when X = 44 AND Y = 128 else
"100010011101" when X = 45 AND Y = 128 else
"100010011101" when X = 46 AND Y = 128 else
"100010011101" when X = 47 AND Y = 128 else
"100010011101" when X = 48 AND Y = 128 else
"100010011101" when X = 49 AND Y = 128 else
"100010011101" when X = 50 AND Y = 128 else
"100010011101" when X = 51 AND Y = 128 else
"100010011101" when X = 52 AND Y = 128 else
"100010011101" when X = 53 AND Y = 128 else
"100010011101" when X = 54 AND Y = 128 else
"100010011101" when X = 55 AND Y = 128 else
"100010011101" when X = 56 AND Y = 128 else
"100010011101" when X = 57 AND Y = 128 else
"100010011101" when X = 58 AND Y = 128 else
"100010011101" when X = 59 AND Y = 128 else
"100010011101" when X = 60 AND Y = 128 else
"100010011101" when X = 61 AND Y = 128 else
"100010011101" when X = 62 AND Y = 128 else
"100010011101" when X = 63 AND Y = 128 else
"100010011101" when X = 64 AND Y = 128 else
"100010011101" when X = 65 AND Y = 128 else
"100010011101" when X = 66 AND Y = 128 else
"100010011101" when X = 67 AND Y = 128 else
"100010011101" when X = 68 AND Y = 128 else
"100010011101" when X = 69 AND Y = 128 else
"100010011101" when X = 70 AND Y = 128 else
"100010011101" when X = 71 AND Y = 128 else
"100010011101" when X = 72 AND Y = 128 else
"100010011101" when X = 73 AND Y = 128 else
"100010011101" when X = 74 AND Y = 128 else
"100010011101" when X = 75 AND Y = 128 else
"100010011101" when X = 76 AND Y = 128 else
"100010011101" when X = 77 AND Y = 128 else
"100010011101" when X = 78 AND Y = 128 else
"100010011101" when X = 79 AND Y = 128 else
"100010011101" when X = 80 AND Y = 128 else
"100010011101" when X = 81 AND Y = 128 else
"100010011101" when X = 82 AND Y = 128 else
"100010011101" when X = 83 AND Y = 128 else
"100010011101" when X = 84 AND Y = 128 else
"100010011101" when X = 85 AND Y = 128 else
"100010011101" when X = 86 AND Y = 128 else
"100010011101" when X = 87 AND Y = 128 else
"100010011101" when X = 88 AND Y = 128 else
"100010011101" when X = 89 AND Y = 128 else
"100010011101" when X = 90 AND Y = 128 else
"100010011101" when X = 91 AND Y = 128 else
"100010011101" when X = 92 AND Y = 128 else
"100010011101" when X = 93 AND Y = 128 else
"100010011101" when X = 94 AND Y = 128 else
"100010011101" when X = 95 AND Y = 128 else
"100010011101" when X = 96 AND Y = 128 else
"100010011101" when X = 97 AND Y = 128 else
"100010011101" when X = 98 AND Y = 128 else
"100010011101" when X = 99 AND Y = 128 else
"100010011101" when X = 100 AND Y = 128 else
"100010011101" when X = 101 AND Y = 128 else
"100010011101" when X = 102 AND Y = 128 else
"100010011101" when X = 103 AND Y = 128 else
"100010011101" when X = 104 AND Y = 128 else
"100010011101" when X = 105 AND Y = 128 else
"100010011101" when X = 106 AND Y = 128 else
"100010011101" when X = 107 AND Y = 128 else
"100010011101" when X = 108 AND Y = 128 else
"100010011101" when X = 109 AND Y = 128 else
"110111011111" when X = 110 AND Y = 128 else
"110111011111" when X = 111 AND Y = 128 else
"110111011111" when X = 112 AND Y = 128 else
"110111011111" when X = 113 AND Y = 128 else
"110111011111" when X = 114 AND Y = 128 else
"110111011111" when X = 115 AND Y = 128 else
"110111011111" when X = 116 AND Y = 128 else
"110111011111" when X = 117 AND Y = 128 else
"110111011111" when X = 118 AND Y = 128 else
"110111011111" when X = 119 AND Y = 128 else
"110111011111" when X = 120 AND Y = 128 else
"110111011111" when X = 121 AND Y = 128 else
"110111011111" when X = 122 AND Y = 128 else
"110111011111" when X = 123 AND Y = 128 else
"110111011111" when X = 124 AND Y = 128 else
"110111011111" when X = 125 AND Y = 128 else
"110111011111" when X = 126 AND Y = 128 else
"110111011111" when X = 127 AND Y = 128 else
"110111011111" when X = 128 AND Y = 128 else
"110111011111" when X = 129 AND Y = 128 else
"110111011111" when X = 130 AND Y = 128 else
"110111011111" when X = 131 AND Y = 128 else
"110111011111" when X = 132 AND Y = 128 else
"110111011111" when X = 133 AND Y = 128 else
"110111011111" when X = 134 AND Y = 128 else
"110111011111" when X = 135 AND Y = 128 else
"110111011111" when X = 136 AND Y = 128 else
"110111011111" when X = 137 AND Y = 128 else
"110111011111" when X = 138 AND Y = 128 else
"110111011111" when X = 139 AND Y = 128 else
"110111011111" when X = 140 AND Y = 128 else
"110111011111" when X = 141 AND Y = 128 else
"110111011111" when X = 142 AND Y = 128 else
"110111011111" when X = 143 AND Y = 128 else
"110111011111" when X = 144 AND Y = 128 else
"110111011111" when X = 145 AND Y = 128 else
"110111011111" when X = 146 AND Y = 128 else
"110111011111" when X = 147 AND Y = 128 else
"110111011111" when X = 148 AND Y = 128 else
"110111011111" when X = 149 AND Y = 128 else
"110111011111" when X = 150 AND Y = 128 else
"110111011111" when X = 151 AND Y = 128 else
"110111011111" when X = 152 AND Y = 128 else
"110111011111" when X = 153 AND Y = 128 else
"110111011111" when X = 154 AND Y = 128 else
"110111011111" when X = 155 AND Y = 128 else
"110111011111" when X = 156 AND Y = 128 else
"110111011111" when X = 157 AND Y = 128 else
"110111011111" when X = 158 AND Y = 128 else
"110111011111" when X = 159 AND Y = 128 else
"110111011111" when X = 160 AND Y = 128 else
"110111011111" when X = 161 AND Y = 128 else
"110111011111" when X = 162 AND Y = 128 else
"110111011111" when X = 163 AND Y = 128 else
"110111011111" when X = 164 AND Y = 128 else
"110111011111" when X = 165 AND Y = 128 else
"110111011111" when X = 166 AND Y = 128 else
"110111011111" when X = 167 AND Y = 128 else
"110111011111" when X = 168 AND Y = 128 else
"110111011111" when X = 169 AND Y = 128 else
"110111011111" when X = 170 AND Y = 128 else
"110111011111" when X = 171 AND Y = 128 else
"110111011111" when X = 172 AND Y = 128 else
"110111011111" when X = 173 AND Y = 128 else
"110111011111" when X = 174 AND Y = 128 else
"110111011111" when X = 175 AND Y = 128 else
"110111011111" when X = 176 AND Y = 128 else
"110111011111" when X = 177 AND Y = 128 else
"110111011111" when X = 178 AND Y = 128 else
"110111011111" when X = 179 AND Y = 128 else
"110111011111" when X = 180 AND Y = 128 else
"110111011111" when X = 181 AND Y = 128 else
"110111011111" when X = 182 AND Y = 128 else
"110111011111" when X = 183 AND Y = 128 else
"110111011111" when X = 184 AND Y = 128 else
"110111011111" when X = 185 AND Y = 128 else
"110111011111" when X = 186 AND Y = 128 else
"110111011111" when X = 187 AND Y = 128 else
"110111011111" when X = 188 AND Y = 128 else
"110111011111" when X = 189 AND Y = 128 else
"110111011111" when X = 190 AND Y = 128 else
"110111011111" when X = 191 AND Y = 128 else
"110111011111" when X = 192 AND Y = 128 else
"110111011111" when X = 193 AND Y = 128 else
"110111011111" when X = 194 AND Y = 128 else
"110111011111" when X = 195 AND Y = 128 else
"110111011111" when X = 196 AND Y = 128 else
"110111011111" when X = 197 AND Y = 128 else
"110111011111" when X = 198 AND Y = 128 else
"110111011111" when X = 199 AND Y = 128 else
"110111011111" when X = 200 AND Y = 128 else
"110111011111" when X = 201 AND Y = 128 else
"110111011111" when X = 202 AND Y = 128 else
"110111011111" when X = 203 AND Y = 128 else
"110111011111" when X = 204 AND Y = 128 else
"110111011111" when X = 205 AND Y = 128 else
"110111011111" when X = 206 AND Y = 128 else
"110111011111" when X = 207 AND Y = 128 else
"110111011111" when X = 208 AND Y = 128 else
"110111011111" when X = 209 AND Y = 128 else
"110111011111" when X = 210 AND Y = 128 else
"110111011111" when X = 211 AND Y = 128 else
"110111011111" when X = 212 AND Y = 128 else
"110111011111" when X = 213 AND Y = 128 else
"110111011111" when X = 214 AND Y = 128 else
"110111011111" when X = 215 AND Y = 128 else
"110111011111" when X = 216 AND Y = 128 else
"110111011111" when X = 217 AND Y = 128 else
"110111011111" when X = 218 AND Y = 128 else
"110111011111" when X = 219 AND Y = 128 else
"110111011111" when X = 220 AND Y = 128 else
"110111011111" when X = 221 AND Y = 128 else
"110111011111" when X = 222 AND Y = 128 else
"110111011111" when X = 223 AND Y = 128 else
"110111011111" when X = 224 AND Y = 128 else
"110111011111" when X = 225 AND Y = 128 else
"110111011111" when X = 226 AND Y = 128 else
"110111011111" when X = 227 AND Y = 128 else
"110111011111" when X = 228 AND Y = 128 else
"110111011111" when X = 229 AND Y = 128 else
"110111011111" when X = 230 AND Y = 128 else
"110111011111" when X = 231 AND Y = 128 else
"110111011111" when X = 232 AND Y = 128 else
"110111011111" when X = 233 AND Y = 128 else
"110111011111" when X = 234 AND Y = 128 else
"000000000000" when X = 235 AND Y = 128 else
"000000000000" when X = 236 AND Y = 128 else
"000000000000" when X = 237 AND Y = 128 else
"000000000000" when X = 238 AND Y = 128 else
"000000000000" when X = 239 AND Y = 128 else
"000000000000" when X = 240 AND Y = 128 else
"000000000000" when X = 241 AND Y = 128 else
"000000000000" when X = 242 AND Y = 128 else
"000000000000" when X = 243 AND Y = 128 else
"000000000000" when X = 244 AND Y = 128 else
"110111011111" when X = 245 AND Y = 128 else
"110111011111" when X = 246 AND Y = 128 else
"110111011111" when X = 247 AND Y = 128 else
"110111011111" when X = 248 AND Y = 128 else
"110111011111" when X = 249 AND Y = 128 else
"110111011111" when X = 250 AND Y = 128 else
"110111011111" when X = 251 AND Y = 128 else
"110111011111" when X = 252 AND Y = 128 else
"110111011111" when X = 253 AND Y = 128 else
"110111011111" when X = 254 AND Y = 128 else
"110111011111" when X = 255 AND Y = 128 else
"110111011111" when X = 256 AND Y = 128 else
"110111011111" when X = 257 AND Y = 128 else
"110111011111" when X = 258 AND Y = 128 else
"110111011111" when X = 259 AND Y = 128 else
"110111011111" when X = 260 AND Y = 128 else
"110111011111" when X = 261 AND Y = 128 else
"110111011111" when X = 262 AND Y = 128 else
"110111011111" when X = 263 AND Y = 128 else
"110111011111" when X = 264 AND Y = 128 else
"110111011111" when X = 265 AND Y = 128 else
"110111011111" when X = 266 AND Y = 128 else
"110111011111" when X = 267 AND Y = 128 else
"110111011111" when X = 268 AND Y = 128 else
"110111011111" when X = 269 AND Y = 128 else
"110111011111" when X = 270 AND Y = 128 else
"110111011111" when X = 271 AND Y = 128 else
"110111011111" when X = 272 AND Y = 128 else
"110111011111" when X = 273 AND Y = 128 else
"110111011111" when X = 274 AND Y = 128 else
"110111011111" when X = 275 AND Y = 128 else
"110111011111" when X = 276 AND Y = 128 else
"110111011111" when X = 277 AND Y = 128 else
"110111011111" when X = 278 AND Y = 128 else
"110111011111" when X = 279 AND Y = 128 else
"110111011111" when X = 280 AND Y = 128 else
"110111011111" when X = 281 AND Y = 128 else
"110111011111" when X = 282 AND Y = 128 else
"110111011111" when X = 283 AND Y = 128 else
"110111011111" when X = 284 AND Y = 128 else
"110111011111" when X = 285 AND Y = 128 else
"110111011111" when X = 286 AND Y = 128 else
"110111011111" when X = 287 AND Y = 128 else
"110111011111" when X = 288 AND Y = 128 else
"110111011111" when X = 289 AND Y = 128 else
"110111011111" when X = 290 AND Y = 128 else
"110111011111" when X = 291 AND Y = 128 else
"110111011111" when X = 292 AND Y = 128 else
"110111011111" when X = 293 AND Y = 128 else
"110111011111" when X = 294 AND Y = 128 else
"110111011111" when X = 295 AND Y = 128 else
"110111011111" when X = 296 AND Y = 128 else
"110111011111" when X = 297 AND Y = 128 else
"110111011111" when X = 298 AND Y = 128 else
"110111011111" when X = 299 AND Y = 128 else
"110111011111" when X = 300 AND Y = 128 else
"110111011111" when X = 301 AND Y = 128 else
"110111011111" when X = 302 AND Y = 128 else
"110111011111" when X = 303 AND Y = 128 else
"110111011111" when X = 304 AND Y = 128 else
"110111011111" when X = 305 AND Y = 128 else
"110111011111" when X = 306 AND Y = 128 else
"110111011111" when X = 307 AND Y = 128 else
"110111011111" when X = 308 AND Y = 128 else
"110111011111" when X = 309 AND Y = 128 else
"110111011111" when X = 310 AND Y = 128 else
"110111011111" when X = 311 AND Y = 128 else
"110111011111" when X = 312 AND Y = 128 else
"110111011111" when X = 313 AND Y = 128 else
"110111011111" when X = 314 AND Y = 128 else
"110111011111" when X = 315 AND Y = 128 else
"110111011111" when X = 316 AND Y = 128 else
"110111011111" when X = 317 AND Y = 128 else
"110111011111" when X = 318 AND Y = 128 else
"110111011111" when X = 319 AND Y = 128 else
"000000000000" when X = 320 AND Y = 128 else
"000000000000" when X = 321 AND Y = 128 else
"000000000000" when X = 322 AND Y = 128 else
"000000000000" when X = 323 AND Y = 128 else
"000000000000" when X = 324 AND Y = 128 else
"100010011101" when X = 0 AND Y = 129 else
"100010011101" when X = 1 AND Y = 129 else
"100010011101" when X = 2 AND Y = 129 else
"100010011101" when X = 3 AND Y = 129 else
"100010011101" when X = 4 AND Y = 129 else
"100010011101" when X = 5 AND Y = 129 else
"100010011101" when X = 6 AND Y = 129 else
"100010011101" when X = 7 AND Y = 129 else
"100010011101" when X = 8 AND Y = 129 else
"100010011101" when X = 9 AND Y = 129 else
"100010011101" when X = 10 AND Y = 129 else
"100010011101" when X = 11 AND Y = 129 else
"100010011101" when X = 12 AND Y = 129 else
"100010011101" when X = 13 AND Y = 129 else
"100010011101" when X = 14 AND Y = 129 else
"100010011101" when X = 15 AND Y = 129 else
"100010011101" when X = 16 AND Y = 129 else
"100010011101" when X = 17 AND Y = 129 else
"100010011101" when X = 18 AND Y = 129 else
"100010011101" when X = 19 AND Y = 129 else
"100010011101" when X = 20 AND Y = 129 else
"100010011101" when X = 21 AND Y = 129 else
"100010011101" when X = 22 AND Y = 129 else
"100010011101" when X = 23 AND Y = 129 else
"100010011101" when X = 24 AND Y = 129 else
"100010011101" when X = 25 AND Y = 129 else
"100010011101" when X = 26 AND Y = 129 else
"100010011101" when X = 27 AND Y = 129 else
"100010011101" when X = 28 AND Y = 129 else
"100010011101" when X = 29 AND Y = 129 else
"100010011101" when X = 30 AND Y = 129 else
"100010011101" when X = 31 AND Y = 129 else
"100010011101" when X = 32 AND Y = 129 else
"100010011101" when X = 33 AND Y = 129 else
"100010011101" when X = 34 AND Y = 129 else
"100010011101" when X = 35 AND Y = 129 else
"100010011101" when X = 36 AND Y = 129 else
"100010011101" when X = 37 AND Y = 129 else
"100010011101" when X = 38 AND Y = 129 else
"100010011101" when X = 39 AND Y = 129 else
"100010011101" when X = 40 AND Y = 129 else
"100010011101" when X = 41 AND Y = 129 else
"100010011101" when X = 42 AND Y = 129 else
"100010011101" when X = 43 AND Y = 129 else
"100010011101" when X = 44 AND Y = 129 else
"100010011101" when X = 45 AND Y = 129 else
"100010011101" when X = 46 AND Y = 129 else
"100010011101" when X = 47 AND Y = 129 else
"100010011101" when X = 48 AND Y = 129 else
"100010011101" when X = 49 AND Y = 129 else
"100010011101" when X = 50 AND Y = 129 else
"100010011101" when X = 51 AND Y = 129 else
"100010011101" when X = 52 AND Y = 129 else
"100010011101" when X = 53 AND Y = 129 else
"100010011101" when X = 54 AND Y = 129 else
"100010011101" when X = 55 AND Y = 129 else
"100010011101" when X = 56 AND Y = 129 else
"100010011101" when X = 57 AND Y = 129 else
"100010011101" when X = 58 AND Y = 129 else
"100010011101" when X = 59 AND Y = 129 else
"100010011101" when X = 60 AND Y = 129 else
"100010011101" when X = 61 AND Y = 129 else
"100010011101" when X = 62 AND Y = 129 else
"100010011101" when X = 63 AND Y = 129 else
"100010011101" when X = 64 AND Y = 129 else
"100010011101" when X = 65 AND Y = 129 else
"100010011101" when X = 66 AND Y = 129 else
"100010011101" when X = 67 AND Y = 129 else
"100010011101" when X = 68 AND Y = 129 else
"100010011101" when X = 69 AND Y = 129 else
"100010011101" when X = 70 AND Y = 129 else
"100010011101" when X = 71 AND Y = 129 else
"100010011101" when X = 72 AND Y = 129 else
"100010011101" when X = 73 AND Y = 129 else
"100010011101" when X = 74 AND Y = 129 else
"100010011101" when X = 75 AND Y = 129 else
"100010011101" when X = 76 AND Y = 129 else
"100010011101" when X = 77 AND Y = 129 else
"100010011101" when X = 78 AND Y = 129 else
"100010011101" when X = 79 AND Y = 129 else
"100010011101" when X = 80 AND Y = 129 else
"100010011101" when X = 81 AND Y = 129 else
"100010011101" when X = 82 AND Y = 129 else
"100010011101" when X = 83 AND Y = 129 else
"100010011101" when X = 84 AND Y = 129 else
"100010011101" when X = 85 AND Y = 129 else
"100010011101" when X = 86 AND Y = 129 else
"100010011101" when X = 87 AND Y = 129 else
"100010011101" when X = 88 AND Y = 129 else
"100010011101" when X = 89 AND Y = 129 else
"100010011101" when X = 90 AND Y = 129 else
"100010011101" when X = 91 AND Y = 129 else
"100010011101" when X = 92 AND Y = 129 else
"100010011101" when X = 93 AND Y = 129 else
"100010011101" when X = 94 AND Y = 129 else
"100010011101" when X = 95 AND Y = 129 else
"100010011101" when X = 96 AND Y = 129 else
"100010011101" when X = 97 AND Y = 129 else
"100010011101" when X = 98 AND Y = 129 else
"100010011101" when X = 99 AND Y = 129 else
"100010011101" when X = 100 AND Y = 129 else
"100010011101" when X = 101 AND Y = 129 else
"100010011101" when X = 102 AND Y = 129 else
"100010011101" when X = 103 AND Y = 129 else
"100010011101" when X = 104 AND Y = 129 else
"100010011101" when X = 105 AND Y = 129 else
"100010011101" when X = 106 AND Y = 129 else
"100010011101" when X = 107 AND Y = 129 else
"100010011101" when X = 108 AND Y = 129 else
"100010011101" when X = 109 AND Y = 129 else
"110111011111" when X = 110 AND Y = 129 else
"110111011111" when X = 111 AND Y = 129 else
"110111011111" when X = 112 AND Y = 129 else
"110111011111" when X = 113 AND Y = 129 else
"110111011111" when X = 114 AND Y = 129 else
"110111011111" when X = 115 AND Y = 129 else
"110111011111" when X = 116 AND Y = 129 else
"110111011111" when X = 117 AND Y = 129 else
"110111011111" when X = 118 AND Y = 129 else
"110111011111" when X = 119 AND Y = 129 else
"110111011111" when X = 120 AND Y = 129 else
"110111011111" when X = 121 AND Y = 129 else
"110111011111" when X = 122 AND Y = 129 else
"110111011111" when X = 123 AND Y = 129 else
"110111011111" when X = 124 AND Y = 129 else
"110111011111" when X = 125 AND Y = 129 else
"110111011111" when X = 126 AND Y = 129 else
"110111011111" when X = 127 AND Y = 129 else
"110111011111" when X = 128 AND Y = 129 else
"110111011111" when X = 129 AND Y = 129 else
"110111011111" when X = 130 AND Y = 129 else
"110111011111" when X = 131 AND Y = 129 else
"110111011111" when X = 132 AND Y = 129 else
"110111011111" when X = 133 AND Y = 129 else
"110111011111" when X = 134 AND Y = 129 else
"110111011111" when X = 135 AND Y = 129 else
"110111011111" when X = 136 AND Y = 129 else
"110111011111" when X = 137 AND Y = 129 else
"110111011111" when X = 138 AND Y = 129 else
"110111011111" when X = 139 AND Y = 129 else
"110111011111" when X = 140 AND Y = 129 else
"110111011111" when X = 141 AND Y = 129 else
"110111011111" when X = 142 AND Y = 129 else
"110111011111" when X = 143 AND Y = 129 else
"110111011111" when X = 144 AND Y = 129 else
"110111011111" when X = 145 AND Y = 129 else
"110111011111" when X = 146 AND Y = 129 else
"110111011111" when X = 147 AND Y = 129 else
"110111011111" when X = 148 AND Y = 129 else
"110111011111" when X = 149 AND Y = 129 else
"110111011111" when X = 150 AND Y = 129 else
"110111011111" when X = 151 AND Y = 129 else
"110111011111" when X = 152 AND Y = 129 else
"110111011111" when X = 153 AND Y = 129 else
"110111011111" when X = 154 AND Y = 129 else
"110111011111" when X = 155 AND Y = 129 else
"110111011111" when X = 156 AND Y = 129 else
"110111011111" when X = 157 AND Y = 129 else
"110111011111" when X = 158 AND Y = 129 else
"110111011111" when X = 159 AND Y = 129 else
"110111011111" when X = 160 AND Y = 129 else
"110111011111" when X = 161 AND Y = 129 else
"110111011111" when X = 162 AND Y = 129 else
"110111011111" when X = 163 AND Y = 129 else
"110111011111" when X = 164 AND Y = 129 else
"110111011111" when X = 165 AND Y = 129 else
"110111011111" when X = 166 AND Y = 129 else
"110111011111" when X = 167 AND Y = 129 else
"110111011111" when X = 168 AND Y = 129 else
"110111011111" when X = 169 AND Y = 129 else
"110111011111" when X = 170 AND Y = 129 else
"110111011111" when X = 171 AND Y = 129 else
"110111011111" when X = 172 AND Y = 129 else
"110111011111" when X = 173 AND Y = 129 else
"110111011111" when X = 174 AND Y = 129 else
"110111011111" when X = 175 AND Y = 129 else
"110111011111" when X = 176 AND Y = 129 else
"110111011111" when X = 177 AND Y = 129 else
"110111011111" when X = 178 AND Y = 129 else
"110111011111" when X = 179 AND Y = 129 else
"110111011111" when X = 180 AND Y = 129 else
"110111011111" when X = 181 AND Y = 129 else
"110111011111" when X = 182 AND Y = 129 else
"110111011111" when X = 183 AND Y = 129 else
"110111011111" when X = 184 AND Y = 129 else
"110111011111" when X = 185 AND Y = 129 else
"110111011111" when X = 186 AND Y = 129 else
"110111011111" when X = 187 AND Y = 129 else
"110111011111" when X = 188 AND Y = 129 else
"110111011111" when X = 189 AND Y = 129 else
"110111011111" when X = 190 AND Y = 129 else
"110111011111" when X = 191 AND Y = 129 else
"110111011111" when X = 192 AND Y = 129 else
"110111011111" when X = 193 AND Y = 129 else
"110111011111" when X = 194 AND Y = 129 else
"110111011111" when X = 195 AND Y = 129 else
"110111011111" when X = 196 AND Y = 129 else
"110111011111" when X = 197 AND Y = 129 else
"110111011111" when X = 198 AND Y = 129 else
"110111011111" when X = 199 AND Y = 129 else
"110111011111" when X = 200 AND Y = 129 else
"110111011111" when X = 201 AND Y = 129 else
"110111011111" when X = 202 AND Y = 129 else
"110111011111" when X = 203 AND Y = 129 else
"110111011111" when X = 204 AND Y = 129 else
"110111011111" when X = 205 AND Y = 129 else
"110111011111" when X = 206 AND Y = 129 else
"110111011111" when X = 207 AND Y = 129 else
"110111011111" when X = 208 AND Y = 129 else
"110111011111" when X = 209 AND Y = 129 else
"110111011111" when X = 210 AND Y = 129 else
"110111011111" when X = 211 AND Y = 129 else
"110111011111" when X = 212 AND Y = 129 else
"110111011111" when X = 213 AND Y = 129 else
"110111011111" when X = 214 AND Y = 129 else
"110111011111" when X = 215 AND Y = 129 else
"110111011111" when X = 216 AND Y = 129 else
"110111011111" when X = 217 AND Y = 129 else
"110111011111" when X = 218 AND Y = 129 else
"110111011111" when X = 219 AND Y = 129 else
"110111011111" when X = 220 AND Y = 129 else
"110111011111" when X = 221 AND Y = 129 else
"110111011111" when X = 222 AND Y = 129 else
"110111011111" when X = 223 AND Y = 129 else
"110111011111" when X = 224 AND Y = 129 else
"110111011111" when X = 225 AND Y = 129 else
"110111011111" when X = 226 AND Y = 129 else
"110111011111" when X = 227 AND Y = 129 else
"110111011111" when X = 228 AND Y = 129 else
"110111011111" when X = 229 AND Y = 129 else
"110111011111" when X = 230 AND Y = 129 else
"110111011111" when X = 231 AND Y = 129 else
"110111011111" when X = 232 AND Y = 129 else
"110111011111" when X = 233 AND Y = 129 else
"110111011111" when X = 234 AND Y = 129 else
"000000000000" when X = 235 AND Y = 129 else
"000000000000" when X = 236 AND Y = 129 else
"000000000000" when X = 237 AND Y = 129 else
"000000000000" when X = 238 AND Y = 129 else
"000000000000" when X = 239 AND Y = 129 else
"000000000000" when X = 240 AND Y = 129 else
"000000000000" when X = 241 AND Y = 129 else
"000000000000" when X = 242 AND Y = 129 else
"000000000000" when X = 243 AND Y = 129 else
"000000000000" when X = 244 AND Y = 129 else
"110111011111" when X = 245 AND Y = 129 else
"110111011111" when X = 246 AND Y = 129 else
"110111011111" when X = 247 AND Y = 129 else
"110111011111" when X = 248 AND Y = 129 else
"110111011111" when X = 249 AND Y = 129 else
"110111011111" when X = 250 AND Y = 129 else
"110111011111" when X = 251 AND Y = 129 else
"110111011111" when X = 252 AND Y = 129 else
"110111011111" when X = 253 AND Y = 129 else
"110111011111" when X = 254 AND Y = 129 else
"110111011111" when X = 255 AND Y = 129 else
"110111011111" when X = 256 AND Y = 129 else
"110111011111" when X = 257 AND Y = 129 else
"110111011111" when X = 258 AND Y = 129 else
"110111011111" when X = 259 AND Y = 129 else
"110111011111" when X = 260 AND Y = 129 else
"110111011111" when X = 261 AND Y = 129 else
"110111011111" when X = 262 AND Y = 129 else
"110111011111" when X = 263 AND Y = 129 else
"110111011111" when X = 264 AND Y = 129 else
"110111011111" when X = 265 AND Y = 129 else
"110111011111" when X = 266 AND Y = 129 else
"110111011111" when X = 267 AND Y = 129 else
"110111011111" when X = 268 AND Y = 129 else
"110111011111" when X = 269 AND Y = 129 else
"110111011111" when X = 270 AND Y = 129 else
"110111011111" when X = 271 AND Y = 129 else
"110111011111" when X = 272 AND Y = 129 else
"110111011111" when X = 273 AND Y = 129 else
"110111011111" when X = 274 AND Y = 129 else
"110111011111" when X = 275 AND Y = 129 else
"110111011111" when X = 276 AND Y = 129 else
"110111011111" when X = 277 AND Y = 129 else
"110111011111" when X = 278 AND Y = 129 else
"110111011111" when X = 279 AND Y = 129 else
"110111011111" when X = 280 AND Y = 129 else
"110111011111" when X = 281 AND Y = 129 else
"110111011111" when X = 282 AND Y = 129 else
"110111011111" when X = 283 AND Y = 129 else
"110111011111" when X = 284 AND Y = 129 else
"110111011111" when X = 285 AND Y = 129 else
"110111011111" when X = 286 AND Y = 129 else
"110111011111" when X = 287 AND Y = 129 else
"110111011111" when X = 288 AND Y = 129 else
"110111011111" when X = 289 AND Y = 129 else
"110111011111" when X = 290 AND Y = 129 else
"110111011111" when X = 291 AND Y = 129 else
"110111011111" when X = 292 AND Y = 129 else
"110111011111" when X = 293 AND Y = 129 else
"110111011111" when X = 294 AND Y = 129 else
"110111011111" when X = 295 AND Y = 129 else
"110111011111" when X = 296 AND Y = 129 else
"110111011111" when X = 297 AND Y = 129 else
"110111011111" when X = 298 AND Y = 129 else
"110111011111" when X = 299 AND Y = 129 else
"110111011111" when X = 300 AND Y = 129 else
"110111011111" when X = 301 AND Y = 129 else
"110111011111" when X = 302 AND Y = 129 else
"110111011111" when X = 303 AND Y = 129 else
"110111011111" when X = 304 AND Y = 129 else
"110111011111" when X = 305 AND Y = 129 else
"110111011111" when X = 306 AND Y = 129 else
"110111011111" when X = 307 AND Y = 129 else
"110111011111" when X = 308 AND Y = 129 else
"110111011111" when X = 309 AND Y = 129 else
"110111011111" when X = 310 AND Y = 129 else
"110111011111" when X = 311 AND Y = 129 else
"110111011111" when X = 312 AND Y = 129 else
"110111011111" when X = 313 AND Y = 129 else
"110111011111" when X = 314 AND Y = 129 else
"110111011111" when X = 315 AND Y = 129 else
"110111011111" when X = 316 AND Y = 129 else
"110111011111" when X = 317 AND Y = 129 else
"110111011111" when X = 318 AND Y = 129 else
"110111011111" when X = 319 AND Y = 129 else
"000000000000" when X = 320 AND Y = 129 else
"000000000000" when X = 321 AND Y = 129 else
"000000000000" when X = 322 AND Y = 129 else
"000000000000" when X = 323 AND Y = 129 else
"000000000000" when X = 324 AND Y = 129 else
"000000000000" when X = 0 AND Y = 130 else
"000000000000" when X = 1 AND Y = 130 else
"000000000000" when X = 2 AND Y = 130 else
"000000000000" when X = 3 AND Y = 130 else
"000000000000" when X = 4 AND Y = 130 else
"000000000000" when X = 5 AND Y = 130 else
"000000000000" when X = 6 AND Y = 130 else
"000000000000" when X = 7 AND Y = 130 else
"000000000000" when X = 8 AND Y = 130 else
"000000000000" when X = 9 AND Y = 130 else
"000000000000" when X = 10 AND Y = 130 else
"000000000000" when X = 11 AND Y = 130 else
"000000000000" when X = 12 AND Y = 130 else
"000000000000" when X = 13 AND Y = 130 else
"000000000000" when X = 14 AND Y = 130 else
"000000000000" when X = 15 AND Y = 130 else
"000000000000" when X = 16 AND Y = 130 else
"000000000000" when X = 17 AND Y = 130 else
"000000000000" when X = 18 AND Y = 130 else
"000000000000" when X = 19 AND Y = 130 else
"000000000000" when X = 20 AND Y = 130 else
"000000000000" when X = 21 AND Y = 130 else
"000000000000" when X = 22 AND Y = 130 else
"000000000000" when X = 23 AND Y = 130 else
"000000000000" when X = 24 AND Y = 130 else
"000000000000" when X = 25 AND Y = 130 else
"000000000000" when X = 26 AND Y = 130 else
"000000000000" when X = 27 AND Y = 130 else
"000000000000" when X = 28 AND Y = 130 else
"000000000000" when X = 29 AND Y = 130 else
"000000000000" when X = 30 AND Y = 130 else
"000000000000" when X = 31 AND Y = 130 else
"000000000000" when X = 32 AND Y = 130 else
"000000000000" when X = 33 AND Y = 130 else
"000000000000" when X = 34 AND Y = 130 else
"000000000000" when X = 35 AND Y = 130 else
"000000000000" when X = 36 AND Y = 130 else
"000000000000" when X = 37 AND Y = 130 else
"000000000000" when X = 38 AND Y = 130 else
"000000000000" when X = 39 AND Y = 130 else
"100010011101" when X = 40 AND Y = 130 else
"100010011101" when X = 41 AND Y = 130 else
"100010011101" when X = 42 AND Y = 130 else
"100010011101" when X = 43 AND Y = 130 else
"100010011101" when X = 44 AND Y = 130 else
"100010011101" when X = 45 AND Y = 130 else
"100010011101" when X = 46 AND Y = 130 else
"100010011101" when X = 47 AND Y = 130 else
"100010011101" when X = 48 AND Y = 130 else
"100010011101" when X = 49 AND Y = 130 else
"100010011101" when X = 50 AND Y = 130 else
"100010011101" when X = 51 AND Y = 130 else
"100010011101" when X = 52 AND Y = 130 else
"100010011101" when X = 53 AND Y = 130 else
"100010011101" when X = 54 AND Y = 130 else
"100010011101" when X = 55 AND Y = 130 else
"100010011101" when X = 56 AND Y = 130 else
"100010011101" when X = 57 AND Y = 130 else
"100010011101" when X = 58 AND Y = 130 else
"100010011101" when X = 59 AND Y = 130 else
"100010011101" when X = 60 AND Y = 130 else
"100010011101" when X = 61 AND Y = 130 else
"100010011101" when X = 62 AND Y = 130 else
"100010011101" when X = 63 AND Y = 130 else
"100010011101" when X = 64 AND Y = 130 else
"100010011101" when X = 65 AND Y = 130 else
"100010011101" when X = 66 AND Y = 130 else
"100010011101" when X = 67 AND Y = 130 else
"100010011101" when X = 68 AND Y = 130 else
"100010011101" when X = 69 AND Y = 130 else
"100010011101" when X = 70 AND Y = 130 else
"100010011101" when X = 71 AND Y = 130 else
"100010011101" when X = 72 AND Y = 130 else
"100010011101" when X = 73 AND Y = 130 else
"100010011101" when X = 74 AND Y = 130 else
"100010011101" when X = 75 AND Y = 130 else
"100010011101" when X = 76 AND Y = 130 else
"100010011101" when X = 77 AND Y = 130 else
"100010011101" when X = 78 AND Y = 130 else
"100010011101" when X = 79 AND Y = 130 else
"100010011101" when X = 80 AND Y = 130 else
"100010011101" when X = 81 AND Y = 130 else
"100010011101" when X = 82 AND Y = 130 else
"100010011101" when X = 83 AND Y = 130 else
"100010011101" when X = 84 AND Y = 130 else
"100010011101" when X = 85 AND Y = 130 else
"100010011101" when X = 86 AND Y = 130 else
"100010011101" when X = 87 AND Y = 130 else
"100010011101" when X = 88 AND Y = 130 else
"100010011101" when X = 89 AND Y = 130 else
"100010011101" when X = 90 AND Y = 130 else
"100010011101" when X = 91 AND Y = 130 else
"100010011101" when X = 92 AND Y = 130 else
"100010011101" when X = 93 AND Y = 130 else
"100010011101" when X = 94 AND Y = 130 else
"100010011101" when X = 95 AND Y = 130 else
"100010011101" when X = 96 AND Y = 130 else
"100010011101" when X = 97 AND Y = 130 else
"100010011101" when X = 98 AND Y = 130 else
"100010011101" when X = 99 AND Y = 130 else
"100010011101" when X = 100 AND Y = 130 else
"100010011101" when X = 101 AND Y = 130 else
"100010011101" when X = 102 AND Y = 130 else
"100010011101" when X = 103 AND Y = 130 else
"100010011101" when X = 104 AND Y = 130 else
"100010011101" when X = 105 AND Y = 130 else
"100010011101" when X = 106 AND Y = 130 else
"100010011101" when X = 107 AND Y = 130 else
"100010011101" when X = 108 AND Y = 130 else
"100010011101" when X = 109 AND Y = 130 else
"110111011111" when X = 110 AND Y = 130 else
"110111011111" when X = 111 AND Y = 130 else
"110111011111" when X = 112 AND Y = 130 else
"110111011111" when X = 113 AND Y = 130 else
"110111011111" when X = 114 AND Y = 130 else
"110111011111" when X = 115 AND Y = 130 else
"110111011111" when X = 116 AND Y = 130 else
"110111011111" when X = 117 AND Y = 130 else
"110111011111" when X = 118 AND Y = 130 else
"110111011111" when X = 119 AND Y = 130 else
"110111011111" when X = 120 AND Y = 130 else
"110111011111" when X = 121 AND Y = 130 else
"110111011111" when X = 122 AND Y = 130 else
"110111011111" when X = 123 AND Y = 130 else
"110111011111" when X = 124 AND Y = 130 else
"110111011111" when X = 125 AND Y = 130 else
"110111011111" when X = 126 AND Y = 130 else
"110111011111" when X = 127 AND Y = 130 else
"110111011111" when X = 128 AND Y = 130 else
"110111011111" when X = 129 AND Y = 130 else
"110111011111" when X = 130 AND Y = 130 else
"110111011111" when X = 131 AND Y = 130 else
"110111011111" when X = 132 AND Y = 130 else
"110111011111" when X = 133 AND Y = 130 else
"110111011111" when X = 134 AND Y = 130 else
"110111011111" when X = 135 AND Y = 130 else
"110111011111" when X = 136 AND Y = 130 else
"110111011111" when X = 137 AND Y = 130 else
"110111011111" when X = 138 AND Y = 130 else
"110111011111" when X = 139 AND Y = 130 else
"110111011111" when X = 140 AND Y = 130 else
"110111011111" when X = 141 AND Y = 130 else
"110111011111" when X = 142 AND Y = 130 else
"110111011111" when X = 143 AND Y = 130 else
"110111011111" when X = 144 AND Y = 130 else
"110111011111" when X = 145 AND Y = 130 else
"110111011111" when X = 146 AND Y = 130 else
"110111011111" when X = 147 AND Y = 130 else
"110111011111" when X = 148 AND Y = 130 else
"110111011111" when X = 149 AND Y = 130 else
"110111011111" when X = 150 AND Y = 130 else
"110111011111" when X = 151 AND Y = 130 else
"110111011111" when X = 152 AND Y = 130 else
"110111011111" when X = 153 AND Y = 130 else
"110111011111" when X = 154 AND Y = 130 else
"110111011111" when X = 155 AND Y = 130 else
"110111011111" when X = 156 AND Y = 130 else
"110111011111" when X = 157 AND Y = 130 else
"110111011111" when X = 158 AND Y = 130 else
"110111011111" when X = 159 AND Y = 130 else
"110111011111" when X = 160 AND Y = 130 else
"110111011111" when X = 161 AND Y = 130 else
"110111011111" when X = 162 AND Y = 130 else
"110111011111" when X = 163 AND Y = 130 else
"110111011111" when X = 164 AND Y = 130 else
"110111011111" when X = 165 AND Y = 130 else
"110111011111" when X = 166 AND Y = 130 else
"110111011111" when X = 167 AND Y = 130 else
"110111011111" when X = 168 AND Y = 130 else
"110111011111" when X = 169 AND Y = 130 else
"110111011111" when X = 170 AND Y = 130 else
"110111011111" when X = 171 AND Y = 130 else
"110111011111" when X = 172 AND Y = 130 else
"110111011111" when X = 173 AND Y = 130 else
"110111011111" when X = 174 AND Y = 130 else
"110111011111" when X = 175 AND Y = 130 else
"110111011111" when X = 176 AND Y = 130 else
"110111011111" when X = 177 AND Y = 130 else
"110111011111" when X = 178 AND Y = 130 else
"110111011111" when X = 179 AND Y = 130 else
"110111011111" when X = 180 AND Y = 130 else
"110111011111" when X = 181 AND Y = 130 else
"110111011111" when X = 182 AND Y = 130 else
"110111011111" when X = 183 AND Y = 130 else
"110111011111" when X = 184 AND Y = 130 else
"110111011111" when X = 185 AND Y = 130 else
"110111011111" when X = 186 AND Y = 130 else
"110111011111" when X = 187 AND Y = 130 else
"110111011111" when X = 188 AND Y = 130 else
"110111011111" when X = 189 AND Y = 130 else
"110111011111" when X = 190 AND Y = 130 else
"110111011111" when X = 191 AND Y = 130 else
"110111011111" when X = 192 AND Y = 130 else
"110111011111" when X = 193 AND Y = 130 else
"110111011111" when X = 194 AND Y = 130 else
"110111011111" when X = 195 AND Y = 130 else
"110111011111" when X = 196 AND Y = 130 else
"110111011111" when X = 197 AND Y = 130 else
"110111011111" when X = 198 AND Y = 130 else
"110111011111" when X = 199 AND Y = 130 else
"000000000000" when X = 200 AND Y = 130 else
"000000000000" when X = 201 AND Y = 130 else
"000000000000" when X = 202 AND Y = 130 else
"000000000000" when X = 203 AND Y = 130 else
"000000000000" when X = 204 AND Y = 130 else
"000000000000" when X = 205 AND Y = 130 else
"000000000000" when X = 206 AND Y = 130 else
"000000000000" when X = 207 AND Y = 130 else
"000000000000" when X = 208 AND Y = 130 else
"000000000000" when X = 209 AND Y = 130 else
"000000000000" when X = 210 AND Y = 130 else
"000000000000" when X = 211 AND Y = 130 else
"000000000000" when X = 212 AND Y = 130 else
"000000000000" when X = 213 AND Y = 130 else
"000000000000" when X = 214 AND Y = 130 else
"000000000000" when X = 215 AND Y = 130 else
"000000000000" when X = 216 AND Y = 130 else
"000000000000" when X = 217 AND Y = 130 else
"000000000000" when X = 218 AND Y = 130 else
"000000000000" when X = 219 AND Y = 130 else
"000000000000" when X = 220 AND Y = 130 else
"000000000000" when X = 221 AND Y = 130 else
"000000000000" when X = 222 AND Y = 130 else
"000000000000" when X = 223 AND Y = 130 else
"000000000000" when X = 224 AND Y = 130 else
"000000000000" when X = 225 AND Y = 130 else
"000000000000" when X = 226 AND Y = 130 else
"000000000000" when X = 227 AND Y = 130 else
"000000000000" when X = 228 AND Y = 130 else
"000000000000" when X = 229 AND Y = 130 else
"000000000000" when X = 230 AND Y = 130 else
"000000000000" when X = 231 AND Y = 130 else
"000000000000" when X = 232 AND Y = 130 else
"000000000000" when X = 233 AND Y = 130 else
"000000000000" when X = 234 AND Y = 130 else
"000000000000" when X = 235 AND Y = 130 else
"000000000000" when X = 236 AND Y = 130 else
"000000000000" when X = 237 AND Y = 130 else
"000000000000" when X = 238 AND Y = 130 else
"000000000000" when X = 239 AND Y = 130 else
"000000000000" when X = 240 AND Y = 130 else
"000000000000" when X = 241 AND Y = 130 else
"000000000000" when X = 242 AND Y = 130 else
"000000000000" when X = 243 AND Y = 130 else
"000000000000" when X = 244 AND Y = 130 else
"000000000000" when X = 245 AND Y = 130 else
"000000000000" when X = 246 AND Y = 130 else
"000000000000" when X = 247 AND Y = 130 else
"000000000000" when X = 248 AND Y = 130 else
"000000000000" when X = 249 AND Y = 130 else
"000000000000" when X = 250 AND Y = 130 else
"000000000000" when X = 251 AND Y = 130 else
"000000000000" when X = 252 AND Y = 130 else
"000000000000" when X = 253 AND Y = 130 else
"000000000000" when X = 254 AND Y = 130 else
"000000000000" when X = 255 AND Y = 130 else
"000000000000" when X = 256 AND Y = 130 else
"000000000000" when X = 257 AND Y = 130 else
"000000000000" when X = 258 AND Y = 130 else
"000000000000" when X = 259 AND Y = 130 else
"000000000000" when X = 260 AND Y = 130 else
"000000000000" when X = 261 AND Y = 130 else
"000000000000" when X = 262 AND Y = 130 else
"000000000000" when X = 263 AND Y = 130 else
"000000000000" when X = 264 AND Y = 130 else
"000000000000" when X = 265 AND Y = 130 else
"000000000000" when X = 266 AND Y = 130 else
"000000000000" when X = 267 AND Y = 130 else
"000000000000" when X = 268 AND Y = 130 else
"000000000000" when X = 269 AND Y = 130 else
"000000000000" when X = 270 AND Y = 130 else
"000000000000" when X = 271 AND Y = 130 else
"000000000000" when X = 272 AND Y = 130 else
"000000000000" when X = 273 AND Y = 130 else
"000000000000" when X = 274 AND Y = 130 else
"000000000000" when X = 275 AND Y = 130 else
"000000000000" when X = 276 AND Y = 130 else
"000000000000" when X = 277 AND Y = 130 else
"000000000000" when X = 278 AND Y = 130 else
"000000000000" when X = 279 AND Y = 130 else
"000000000000" when X = 280 AND Y = 130 else
"000000000000" when X = 281 AND Y = 130 else
"000000000000" when X = 282 AND Y = 130 else
"000000000000" when X = 283 AND Y = 130 else
"000000000000" when X = 284 AND Y = 130 else
"000000000000" when X = 285 AND Y = 130 else
"000000000000" when X = 286 AND Y = 130 else
"000000000000" when X = 287 AND Y = 130 else
"000000000000" when X = 288 AND Y = 130 else
"000000000000" when X = 289 AND Y = 130 else
"000000000000" when X = 290 AND Y = 130 else
"000000000000" when X = 291 AND Y = 130 else
"000000000000" when X = 292 AND Y = 130 else
"000000000000" when X = 293 AND Y = 130 else
"000000000000" when X = 294 AND Y = 130 else
"000000000000" when X = 295 AND Y = 130 else
"000000000000" when X = 296 AND Y = 130 else
"000000000000" when X = 297 AND Y = 130 else
"000000000000" when X = 298 AND Y = 130 else
"000000000000" when X = 299 AND Y = 130 else
"000000000000" when X = 300 AND Y = 130 else
"000000000000" when X = 301 AND Y = 130 else
"000000000000" when X = 302 AND Y = 130 else
"000000000000" when X = 303 AND Y = 130 else
"000000000000" when X = 304 AND Y = 130 else
"000000000000" when X = 305 AND Y = 130 else
"000000000000" when X = 306 AND Y = 130 else
"000000000000" when X = 307 AND Y = 130 else
"000000000000" when X = 308 AND Y = 130 else
"000000000000" when X = 309 AND Y = 130 else
"000000000000" when X = 310 AND Y = 130 else
"000000000000" when X = 311 AND Y = 130 else
"000000000000" when X = 312 AND Y = 130 else
"000000000000" when X = 313 AND Y = 130 else
"000000000000" when X = 314 AND Y = 130 else
"000000000000" when X = 315 AND Y = 130 else
"000000000000" when X = 316 AND Y = 130 else
"000000000000" when X = 317 AND Y = 130 else
"000000000000" when X = 318 AND Y = 130 else
"000000000000" when X = 319 AND Y = 130 else
"000000000000" when X = 320 AND Y = 130 else
"000000000000" when X = 321 AND Y = 130 else
"000000000000" when X = 322 AND Y = 130 else
"000000000000" when X = 323 AND Y = 130 else
"000000000000" when X = 324 AND Y = 130 else
"000000000000" when X = 0 AND Y = 131 else
"000000000000" when X = 1 AND Y = 131 else
"000000000000" when X = 2 AND Y = 131 else
"000000000000" when X = 3 AND Y = 131 else
"000000000000" when X = 4 AND Y = 131 else
"000000000000" when X = 5 AND Y = 131 else
"000000000000" when X = 6 AND Y = 131 else
"000000000000" when X = 7 AND Y = 131 else
"000000000000" when X = 8 AND Y = 131 else
"000000000000" when X = 9 AND Y = 131 else
"000000000000" when X = 10 AND Y = 131 else
"000000000000" when X = 11 AND Y = 131 else
"000000000000" when X = 12 AND Y = 131 else
"000000000000" when X = 13 AND Y = 131 else
"000000000000" when X = 14 AND Y = 131 else
"000000000000" when X = 15 AND Y = 131 else
"000000000000" when X = 16 AND Y = 131 else
"000000000000" when X = 17 AND Y = 131 else
"000000000000" when X = 18 AND Y = 131 else
"000000000000" when X = 19 AND Y = 131 else
"000000000000" when X = 20 AND Y = 131 else
"000000000000" when X = 21 AND Y = 131 else
"000000000000" when X = 22 AND Y = 131 else
"000000000000" when X = 23 AND Y = 131 else
"000000000000" when X = 24 AND Y = 131 else
"000000000000" when X = 25 AND Y = 131 else
"000000000000" when X = 26 AND Y = 131 else
"000000000000" when X = 27 AND Y = 131 else
"000000000000" when X = 28 AND Y = 131 else
"000000000000" when X = 29 AND Y = 131 else
"000000000000" when X = 30 AND Y = 131 else
"000000000000" when X = 31 AND Y = 131 else
"000000000000" when X = 32 AND Y = 131 else
"000000000000" when X = 33 AND Y = 131 else
"000000000000" when X = 34 AND Y = 131 else
"000000000000" when X = 35 AND Y = 131 else
"000000000000" when X = 36 AND Y = 131 else
"000000000000" when X = 37 AND Y = 131 else
"000000000000" when X = 38 AND Y = 131 else
"000000000000" when X = 39 AND Y = 131 else
"100010011101" when X = 40 AND Y = 131 else
"100010011101" when X = 41 AND Y = 131 else
"100010011101" when X = 42 AND Y = 131 else
"100010011101" when X = 43 AND Y = 131 else
"100010011101" when X = 44 AND Y = 131 else
"100010011101" when X = 45 AND Y = 131 else
"100010011101" when X = 46 AND Y = 131 else
"100010011101" when X = 47 AND Y = 131 else
"100010011101" when X = 48 AND Y = 131 else
"100010011101" when X = 49 AND Y = 131 else
"100010011101" when X = 50 AND Y = 131 else
"100010011101" when X = 51 AND Y = 131 else
"100010011101" when X = 52 AND Y = 131 else
"100010011101" when X = 53 AND Y = 131 else
"100010011101" when X = 54 AND Y = 131 else
"100010011101" when X = 55 AND Y = 131 else
"100010011101" when X = 56 AND Y = 131 else
"100010011101" when X = 57 AND Y = 131 else
"100010011101" when X = 58 AND Y = 131 else
"100010011101" when X = 59 AND Y = 131 else
"100010011101" when X = 60 AND Y = 131 else
"100010011101" when X = 61 AND Y = 131 else
"100010011101" when X = 62 AND Y = 131 else
"100010011101" when X = 63 AND Y = 131 else
"100010011101" when X = 64 AND Y = 131 else
"100010011101" when X = 65 AND Y = 131 else
"100010011101" when X = 66 AND Y = 131 else
"100010011101" when X = 67 AND Y = 131 else
"100010011101" when X = 68 AND Y = 131 else
"100010011101" when X = 69 AND Y = 131 else
"100010011101" when X = 70 AND Y = 131 else
"100010011101" when X = 71 AND Y = 131 else
"100010011101" when X = 72 AND Y = 131 else
"100010011101" when X = 73 AND Y = 131 else
"100010011101" when X = 74 AND Y = 131 else
"100010011101" when X = 75 AND Y = 131 else
"100010011101" when X = 76 AND Y = 131 else
"100010011101" when X = 77 AND Y = 131 else
"100010011101" when X = 78 AND Y = 131 else
"100010011101" when X = 79 AND Y = 131 else
"100010011101" when X = 80 AND Y = 131 else
"100010011101" when X = 81 AND Y = 131 else
"100010011101" when X = 82 AND Y = 131 else
"100010011101" when X = 83 AND Y = 131 else
"100010011101" when X = 84 AND Y = 131 else
"100010011101" when X = 85 AND Y = 131 else
"100010011101" when X = 86 AND Y = 131 else
"100010011101" when X = 87 AND Y = 131 else
"100010011101" when X = 88 AND Y = 131 else
"100010011101" when X = 89 AND Y = 131 else
"100010011101" when X = 90 AND Y = 131 else
"100010011101" when X = 91 AND Y = 131 else
"100010011101" when X = 92 AND Y = 131 else
"100010011101" when X = 93 AND Y = 131 else
"100010011101" when X = 94 AND Y = 131 else
"100010011101" when X = 95 AND Y = 131 else
"100010011101" when X = 96 AND Y = 131 else
"100010011101" when X = 97 AND Y = 131 else
"100010011101" when X = 98 AND Y = 131 else
"100010011101" when X = 99 AND Y = 131 else
"100010011101" when X = 100 AND Y = 131 else
"100010011101" when X = 101 AND Y = 131 else
"100010011101" when X = 102 AND Y = 131 else
"100010011101" when X = 103 AND Y = 131 else
"100010011101" when X = 104 AND Y = 131 else
"100010011101" when X = 105 AND Y = 131 else
"100010011101" when X = 106 AND Y = 131 else
"100010011101" when X = 107 AND Y = 131 else
"100010011101" when X = 108 AND Y = 131 else
"100010011101" when X = 109 AND Y = 131 else
"110111011111" when X = 110 AND Y = 131 else
"110111011111" when X = 111 AND Y = 131 else
"110111011111" when X = 112 AND Y = 131 else
"110111011111" when X = 113 AND Y = 131 else
"110111011111" when X = 114 AND Y = 131 else
"110111011111" when X = 115 AND Y = 131 else
"110111011111" when X = 116 AND Y = 131 else
"110111011111" when X = 117 AND Y = 131 else
"110111011111" when X = 118 AND Y = 131 else
"110111011111" when X = 119 AND Y = 131 else
"110111011111" when X = 120 AND Y = 131 else
"110111011111" when X = 121 AND Y = 131 else
"110111011111" when X = 122 AND Y = 131 else
"110111011111" when X = 123 AND Y = 131 else
"110111011111" when X = 124 AND Y = 131 else
"110111011111" when X = 125 AND Y = 131 else
"110111011111" when X = 126 AND Y = 131 else
"110111011111" when X = 127 AND Y = 131 else
"110111011111" when X = 128 AND Y = 131 else
"110111011111" when X = 129 AND Y = 131 else
"110111011111" when X = 130 AND Y = 131 else
"110111011111" when X = 131 AND Y = 131 else
"110111011111" when X = 132 AND Y = 131 else
"110111011111" when X = 133 AND Y = 131 else
"110111011111" when X = 134 AND Y = 131 else
"110111011111" when X = 135 AND Y = 131 else
"110111011111" when X = 136 AND Y = 131 else
"110111011111" when X = 137 AND Y = 131 else
"110111011111" when X = 138 AND Y = 131 else
"110111011111" when X = 139 AND Y = 131 else
"110111011111" when X = 140 AND Y = 131 else
"110111011111" when X = 141 AND Y = 131 else
"110111011111" when X = 142 AND Y = 131 else
"110111011111" when X = 143 AND Y = 131 else
"110111011111" when X = 144 AND Y = 131 else
"110111011111" when X = 145 AND Y = 131 else
"110111011111" when X = 146 AND Y = 131 else
"110111011111" when X = 147 AND Y = 131 else
"110111011111" when X = 148 AND Y = 131 else
"110111011111" when X = 149 AND Y = 131 else
"110111011111" when X = 150 AND Y = 131 else
"110111011111" when X = 151 AND Y = 131 else
"110111011111" when X = 152 AND Y = 131 else
"110111011111" when X = 153 AND Y = 131 else
"110111011111" when X = 154 AND Y = 131 else
"110111011111" when X = 155 AND Y = 131 else
"110111011111" when X = 156 AND Y = 131 else
"110111011111" when X = 157 AND Y = 131 else
"110111011111" when X = 158 AND Y = 131 else
"110111011111" when X = 159 AND Y = 131 else
"110111011111" when X = 160 AND Y = 131 else
"110111011111" when X = 161 AND Y = 131 else
"110111011111" when X = 162 AND Y = 131 else
"110111011111" when X = 163 AND Y = 131 else
"110111011111" when X = 164 AND Y = 131 else
"110111011111" when X = 165 AND Y = 131 else
"110111011111" when X = 166 AND Y = 131 else
"110111011111" when X = 167 AND Y = 131 else
"110111011111" when X = 168 AND Y = 131 else
"110111011111" when X = 169 AND Y = 131 else
"110111011111" when X = 170 AND Y = 131 else
"110111011111" when X = 171 AND Y = 131 else
"110111011111" when X = 172 AND Y = 131 else
"110111011111" when X = 173 AND Y = 131 else
"110111011111" when X = 174 AND Y = 131 else
"110111011111" when X = 175 AND Y = 131 else
"110111011111" when X = 176 AND Y = 131 else
"110111011111" when X = 177 AND Y = 131 else
"110111011111" when X = 178 AND Y = 131 else
"110111011111" when X = 179 AND Y = 131 else
"110111011111" when X = 180 AND Y = 131 else
"110111011111" when X = 181 AND Y = 131 else
"110111011111" when X = 182 AND Y = 131 else
"110111011111" when X = 183 AND Y = 131 else
"110111011111" when X = 184 AND Y = 131 else
"110111011111" when X = 185 AND Y = 131 else
"110111011111" when X = 186 AND Y = 131 else
"110111011111" when X = 187 AND Y = 131 else
"110111011111" when X = 188 AND Y = 131 else
"110111011111" when X = 189 AND Y = 131 else
"110111011111" when X = 190 AND Y = 131 else
"110111011111" when X = 191 AND Y = 131 else
"110111011111" when X = 192 AND Y = 131 else
"110111011111" when X = 193 AND Y = 131 else
"110111011111" when X = 194 AND Y = 131 else
"110111011111" when X = 195 AND Y = 131 else
"110111011111" when X = 196 AND Y = 131 else
"110111011111" when X = 197 AND Y = 131 else
"110111011111" when X = 198 AND Y = 131 else
"110111011111" when X = 199 AND Y = 131 else
"000000000000" when X = 200 AND Y = 131 else
"000000000000" when X = 201 AND Y = 131 else
"000000000000" when X = 202 AND Y = 131 else
"000000000000" when X = 203 AND Y = 131 else
"000000000000" when X = 204 AND Y = 131 else
"000000000000" when X = 205 AND Y = 131 else
"000000000000" when X = 206 AND Y = 131 else
"000000000000" when X = 207 AND Y = 131 else
"000000000000" when X = 208 AND Y = 131 else
"000000000000" when X = 209 AND Y = 131 else
"000000000000" when X = 210 AND Y = 131 else
"000000000000" when X = 211 AND Y = 131 else
"000000000000" when X = 212 AND Y = 131 else
"000000000000" when X = 213 AND Y = 131 else
"000000000000" when X = 214 AND Y = 131 else
"000000000000" when X = 215 AND Y = 131 else
"000000000000" when X = 216 AND Y = 131 else
"000000000000" when X = 217 AND Y = 131 else
"000000000000" when X = 218 AND Y = 131 else
"000000000000" when X = 219 AND Y = 131 else
"000000000000" when X = 220 AND Y = 131 else
"000000000000" when X = 221 AND Y = 131 else
"000000000000" when X = 222 AND Y = 131 else
"000000000000" when X = 223 AND Y = 131 else
"000000000000" when X = 224 AND Y = 131 else
"000000000000" when X = 225 AND Y = 131 else
"000000000000" when X = 226 AND Y = 131 else
"000000000000" when X = 227 AND Y = 131 else
"000000000000" when X = 228 AND Y = 131 else
"000000000000" when X = 229 AND Y = 131 else
"000000000000" when X = 230 AND Y = 131 else
"000000000000" when X = 231 AND Y = 131 else
"000000000000" when X = 232 AND Y = 131 else
"000000000000" when X = 233 AND Y = 131 else
"000000000000" when X = 234 AND Y = 131 else
"000000000000" when X = 235 AND Y = 131 else
"000000000000" when X = 236 AND Y = 131 else
"000000000000" when X = 237 AND Y = 131 else
"000000000000" when X = 238 AND Y = 131 else
"000000000000" when X = 239 AND Y = 131 else
"000000000000" when X = 240 AND Y = 131 else
"000000000000" when X = 241 AND Y = 131 else
"000000000000" when X = 242 AND Y = 131 else
"000000000000" when X = 243 AND Y = 131 else
"000000000000" when X = 244 AND Y = 131 else
"000000000000" when X = 245 AND Y = 131 else
"000000000000" when X = 246 AND Y = 131 else
"000000000000" when X = 247 AND Y = 131 else
"000000000000" when X = 248 AND Y = 131 else
"000000000000" when X = 249 AND Y = 131 else
"000000000000" when X = 250 AND Y = 131 else
"000000000000" when X = 251 AND Y = 131 else
"000000000000" when X = 252 AND Y = 131 else
"000000000000" when X = 253 AND Y = 131 else
"000000000000" when X = 254 AND Y = 131 else
"000000000000" when X = 255 AND Y = 131 else
"000000000000" when X = 256 AND Y = 131 else
"000000000000" when X = 257 AND Y = 131 else
"000000000000" when X = 258 AND Y = 131 else
"000000000000" when X = 259 AND Y = 131 else
"000000000000" when X = 260 AND Y = 131 else
"000000000000" when X = 261 AND Y = 131 else
"000000000000" when X = 262 AND Y = 131 else
"000000000000" when X = 263 AND Y = 131 else
"000000000000" when X = 264 AND Y = 131 else
"000000000000" when X = 265 AND Y = 131 else
"000000000000" when X = 266 AND Y = 131 else
"000000000000" when X = 267 AND Y = 131 else
"000000000000" when X = 268 AND Y = 131 else
"000000000000" when X = 269 AND Y = 131 else
"000000000000" when X = 270 AND Y = 131 else
"000000000000" when X = 271 AND Y = 131 else
"000000000000" when X = 272 AND Y = 131 else
"000000000000" when X = 273 AND Y = 131 else
"000000000000" when X = 274 AND Y = 131 else
"000000000000" when X = 275 AND Y = 131 else
"000000000000" when X = 276 AND Y = 131 else
"000000000000" when X = 277 AND Y = 131 else
"000000000000" when X = 278 AND Y = 131 else
"000000000000" when X = 279 AND Y = 131 else
"000000000000" when X = 280 AND Y = 131 else
"000000000000" when X = 281 AND Y = 131 else
"000000000000" when X = 282 AND Y = 131 else
"000000000000" when X = 283 AND Y = 131 else
"000000000000" when X = 284 AND Y = 131 else
"000000000000" when X = 285 AND Y = 131 else
"000000000000" when X = 286 AND Y = 131 else
"000000000000" when X = 287 AND Y = 131 else
"000000000000" when X = 288 AND Y = 131 else
"000000000000" when X = 289 AND Y = 131 else
"000000000000" when X = 290 AND Y = 131 else
"000000000000" when X = 291 AND Y = 131 else
"000000000000" when X = 292 AND Y = 131 else
"000000000000" when X = 293 AND Y = 131 else
"000000000000" when X = 294 AND Y = 131 else
"000000000000" when X = 295 AND Y = 131 else
"000000000000" when X = 296 AND Y = 131 else
"000000000000" when X = 297 AND Y = 131 else
"000000000000" when X = 298 AND Y = 131 else
"000000000000" when X = 299 AND Y = 131 else
"000000000000" when X = 300 AND Y = 131 else
"000000000000" when X = 301 AND Y = 131 else
"000000000000" when X = 302 AND Y = 131 else
"000000000000" when X = 303 AND Y = 131 else
"000000000000" when X = 304 AND Y = 131 else
"000000000000" when X = 305 AND Y = 131 else
"000000000000" when X = 306 AND Y = 131 else
"000000000000" when X = 307 AND Y = 131 else
"000000000000" when X = 308 AND Y = 131 else
"000000000000" when X = 309 AND Y = 131 else
"000000000000" when X = 310 AND Y = 131 else
"000000000000" when X = 311 AND Y = 131 else
"000000000000" when X = 312 AND Y = 131 else
"000000000000" when X = 313 AND Y = 131 else
"000000000000" when X = 314 AND Y = 131 else
"000000000000" when X = 315 AND Y = 131 else
"000000000000" when X = 316 AND Y = 131 else
"000000000000" when X = 317 AND Y = 131 else
"000000000000" when X = 318 AND Y = 131 else
"000000000000" when X = 319 AND Y = 131 else
"000000000000" when X = 320 AND Y = 131 else
"000000000000" when X = 321 AND Y = 131 else
"000000000000" when X = 322 AND Y = 131 else
"000000000000" when X = 323 AND Y = 131 else
"000000000000" when X = 324 AND Y = 131 else
"000000000000" when X = 0 AND Y = 132 else
"000000000000" when X = 1 AND Y = 132 else
"000000000000" when X = 2 AND Y = 132 else
"000000000000" when X = 3 AND Y = 132 else
"000000000000" when X = 4 AND Y = 132 else
"000000000000" when X = 5 AND Y = 132 else
"000000000000" when X = 6 AND Y = 132 else
"000000000000" when X = 7 AND Y = 132 else
"000000000000" when X = 8 AND Y = 132 else
"000000000000" when X = 9 AND Y = 132 else
"000000000000" when X = 10 AND Y = 132 else
"000000000000" when X = 11 AND Y = 132 else
"000000000000" when X = 12 AND Y = 132 else
"000000000000" when X = 13 AND Y = 132 else
"000000000000" when X = 14 AND Y = 132 else
"000000000000" when X = 15 AND Y = 132 else
"000000000000" when X = 16 AND Y = 132 else
"000000000000" when X = 17 AND Y = 132 else
"000000000000" when X = 18 AND Y = 132 else
"000000000000" when X = 19 AND Y = 132 else
"000000000000" when X = 20 AND Y = 132 else
"000000000000" when X = 21 AND Y = 132 else
"000000000000" when X = 22 AND Y = 132 else
"000000000000" when X = 23 AND Y = 132 else
"000000000000" when X = 24 AND Y = 132 else
"000000000000" when X = 25 AND Y = 132 else
"000000000000" when X = 26 AND Y = 132 else
"000000000000" when X = 27 AND Y = 132 else
"000000000000" when X = 28 AND Y = 132 else
"000000000000" when X = 29 AND Y = 132 else
"000000000000" when X = 30 AND Y = 132 else
"000000000000" when X = 31 AND Y = 132 else
"000000000000" when X = 32 AND Y = 132 else
"000000000000" when X = 33 AND Y = 132 else
"000000000000" when X = 34 AND Y = 132 else
"000000000000" when X = 35 AND Y = 132 else
"000000000000" when X = 36 AND Y = 132 else
"000000000000" when X = 37 AND Y = 132 else
"000000000000" when X = 38 AND Y = 132 else
"000000000000" when X = 39 AND Y = 132 else
"100010011101" when X = 40 AND Y = 132 else
"100010011101" when X = 41 AND Y = 132 else
"100010011101" when X = 42 AND Y = 132 else
"100010011101" when X = 43 AND Y = 132 else
"100010011101" when X = 44 AND Y = 132 else
"100010011101" when X = 45 AND Y = 132 else
"100010011101" when X = 46 AND Y = 132 else
"100010011101" when X = 47 AND Y = 132 else
"100010011101" when X = 48 AND Y = 132 else
"100010011101" when X = 49 AND Y = 132 else
"100010011101" when X = 50 AND Y = 132 else
"100010011101" when X = 51 AND Y = 132 else
"100010011101" when X = 52 AND Y = 132 else
"100010011101" when X = 53 AND Y = 132 else
"100010011101" when X = 54 AND Y = 132 else
"100010011101" when X = 55 AND Y = 132 else
"100010011101" when X = 56 AND Y = 132 else
"100010011101" when X = 57 AND Y = 132 else
"100010011101" when X = 58 AND Y = 132 else
"100010011101" when X = 59 AND Y = 132 else
"100010011101" when X = 60 AND Y = 132 else
"100010011101" when X = 61 AND Y = 132 else
"100010011101" when X = 62 AND Y = 132 else
"100010011101" when X = 63 AND Y = 132 else
"100010011101" when X = 64 AND Y = 132 else
"100010011101" when X = 65 AND Y = 132 else
"100010011101" when X = 66 AND Y = 132 else
"100010011101" when X = 67 AND Y = 132 else
"100010011101" when X = 68 AND Y = 132 else
"100010011101" when X = 69 AND Y = 132 else
"100010011101" when X = 70 AND Y = 132 else
"100010011101" when X = 71 AND Y = 132 else
"100010011101" when X = 72 AND Y = 132 else
"100010011101" when X = 73 AND Y = 132 else
"100010011101" when X = 74 AND Y = 132 else
"100010011101" when X = 75 AND Y = 132 else
"100010011101" when X = 76 AND Y = 132 else
"100010011101" when X = 77 AND Y = 132 else
"100010011101" when X = 78 AND Y = 132 else
"100010011101" when X = 79 AND Y = 132 else
"100010011101" when X = 80 AND Y = 132 else
"100010011101" when X = 81 AND Y = 132 else
"100010011101" when X = 82 AND Y = 132 else
"100010011101" when X = 83 AND Y = 132 else
"100010011101" when X = 84 AND Y = 132 else
"100010011101" when X = 85 AND Y = 132 else
"100010011101" when X = 86 AND Y = 132 else
"100010011101" when X = 87 AND Y = 132 else
"100010011101" when X = 88 AND Y = 132 else
"100010011101" when X = 89 AND Y = 132 else
"100010011101" when X = 90 AND Y = 132 else
"100010011101" when X = 91 AND Y = 132 else
"100010011101" when X = 92 AND Y = 132 else
"100010011101" when X = 93 AND Y = 132 else
"100010011101" when X = 94 AND Y = 132 else
"100010011101" when X = 95 AND Y = 132 else
"100010011101" when X = 96 AND Y = 132 else
"100010011101" when X = 97 AND Y = 132 else
"100010011101" when X = 98 AND Y = 132 else
"100010011101" when X = 99 AND Y = 132 else
"100010011101" when X = 100 AND Y = 132 else
"100010011101" when X = 101 AND Y = 132 else
"100010011101" when X = 102 AND Y = 132 else
"100010011101" when X = 103 AND Y = 132 else
"100010011101" when X = 104 AND Y = 132 else
"100010011101" when X = 105 AND Y = 132 else
"100010011101" when X = 106 AND Y = 132 else
"100010011101" when X = 107 AND Y = 132 else
"100010011101" when X = 108 AND Y = 132 else
"100010011101" when X = 109 AND Y = 132 else
"110111011111" when X = 110 AND Y = 132 else
"110111011111" when X = 111 AND Y = 132 else
"110111011111" when X = 112 AND Y = 132 else
"110111011111" when X = 113 AND Y = 132 else
"110111011111" when X = 114 AND Y = 132 else
"110111011111" when X = 115 AND Y = 132 else
"110111011111" when X = 116 AND Y = 132 else
"110111011111" when X = 117 AND Y = 132 else
"110111011111" when X = 118 AND Y = 132 else
"110111011111" when X = 119 AND Y = 132 else
"110111011111" when X = 120 AND Y = 132 else
"110111011111" when X = 121 AND Y = 132 else
"110111011111" when X = 122 AND Y = 132 else
"110111011111" when X = 123 AND Y = 132 else
"110111011111" when X = 124 AND Y = 132 else
"110111011111" when X = 125 AND Y = 132 else
"110111011111" when X = 126 AND Y = 132 else
"110111011111" when X = 127 AND Y = 132 else
"110111011111" when X = 128 AND Y = 132 else
"110111011111" when X = 129 AND Y = 132 else
"110111011111" when X = 130 AND Y = 132 else
"110111011111" when X = 131 AND Y = 132 else
"110111011111" when X = 132 AND Y = 132 else
"110111011111" when X = 133 AND Y = 132 else
"110111011111" when X = 134 AND Y = 132 else
"110111011111" when X = 135 AND Y = 132 else
"110111011111" when X = 136 AND Y = 132 else
"110111011111" when X = 137 AND Y = 132 else
"110111011111" when X = 138 AND Y = 132 else
"110111011111" when X = 139 AND Y = 132 else
"110111011111" when X = 140 AND Y = 132 else
"110111011111" when X = 141 AND Y = 132 else
"110111011111" when X = 142 AND Y = 132 else
"110111011111" when X = 143 AND Y = 132 else
"110111011111" when X = 144 AND Y = 132 else
"110111011111" when X = 145 AND Y = 132 else
"110111011111" when X = 146 AND Y = 132 else
"110111011111" when X = 147 AND Y = 132 else
"110111011111" when X = 148 AND Y = 132 else
"110111011111" when X = 149 AND Y = 132 else
"110111011111" when X = 150 AND Y = 132 else
"110111011111" when X = 151 AND Y = 132 else
"110111011111" when X = 152 AND Y = 132 else
"110111011111" when X = 153 AND Y = 132 else
"110111011111" when X = 154 AND Y = 132 else
"110111011111" when X = 155 AND Y = 132 else
"110111011111" when X = 156 AND Y = 132 else
"110111011111" when X = 157 AND Y = 132 else
"110111011111" when X = 158 AND Y = 132 else
"110111011111" when X = 159 AND Y = 132 else
"110111011111" when X = 160 AND Y = 132 else
"110111011111" when X = 161 AND Y = 132 else
"110111011111" when X = 162 AND Y = 132 else
"110111011111" when X = 163 AND Y = 132 else
"110111011111" when X = 164 AND Y = 132 else
"110111011111" when X = 165 AND Y = 132 else
"110111011111" when X = 166 AND Y = 132 else
"110111011111" when X = 167 AND Y = 132 else
"110111011111" when X = 168 AND Y = 132 else
"110111011111" when X = 169 AND Y = 132 else
"110111011111" when X = 170 AND Y = 132 else
"110111011111" when X = 171 AND Y = 132 else
"110111011111" when X = 172 AND Y = 132 else
"110111011111" when X = 173 AND Y = 132 else
"110111011111" when X = 174 AND Y = 132 else
"110111011111" when X = 175 AND Y = 132 else
"110111011111" when X = 176 AND Y = 132 else
"110111011111" when X = 177 AND Y = 132 else
"110111011111" when X = 178 AND Y = 132 else
"110111011111" when X = 179 AND Y = 132 else
"110111011111" when X = 180 AND Y = 132 else
"110111011111" when X = 181 AND Y = 132 else
"110111011111" when X = 182 AND Y = 132 else
"110111011111" when X = 183 AND Y = 132 else
"110111011111" when X = 184 AND Y = 132 else
"110111011111" when X = 185 AND Y = 132 else
"110111011111" when X = 186 AND Y = 132 else
"110111011111" when X = 187 AND Y = 132 else
"110111011111" when X = 188 AND Y = 132 else
"110111011111" when X = 189 AND Y = 132 else
"110111011111" when X = 190 AND Y = 132 else
"110111011111" when X = 191 AND Y = 132 else
"110111011111" when X = 192 AND Y = 132 else
"110111011111" when X = 193 AND Y = 132 else
"110111011111" when X = 194 AND Y = 132 else
"110111011111" when X = 195 AND Y = 132 else
"110111011111" when X = 196 AND Y = 132 else
"110111011111" when X = 197 AND Y = 132 else
"110111011111" when X = 198 AND Y = 132 else
"110111011111" when X = 199 AND Y = 132 else
"000000000000" when X = 200 AND Y = 132 else
"000000000000" when X = 201 AND Y = 132 else
"000000000000" when X = 202 AND Y = 132 else
"000000000000" when X = 203 AND Y = 132 else
"000000000000" when X = 204 AND Y = 132 else
"000000000000" when X = 205 AND Y = 132 else
"000000000000" when X = 206 AND Y = 132 else
"000000000000" when X = 207 AND Y = 132 else
"000000000000" when X = 208 AND Y = 132 else
"000000000000" when X = 209 AND Y = 132 else
"000000000000" when X = 210 AND Y = 132 else
"000000000000" when X = 211 AND Y = 132 else
"000000000000" when X = 212 AND Y = 132 else
"000000000000" when X = 213 AND Y = 132 else
"000000000000" when X = 214 AND Y = 132 else
"000000000000" when X = 215 AND Y = 132 else
"000000000000" when X = 216 AND Y = 132 else
"000000000000" when X = 217 AND Y = 132 else
"000000000000" when X = 218 AND Y = 132 else
"000000000000" when X = 219 AND Y = 132 else
"000000000000" when X = 220 AND Y = 132 else
"000000000000" when X = 221 AND Y = 132 else
"000000000000" when X = 222 AND Y = 132 else
"000000000000" when X = 223 AND Y = 132 else
"000000000000" when X = 224 AND Y = 132 else
"000000000000" when X = 225 AND Y = 132 else
"000000000000" when X = 226 AND Y = 132 else
"000000000000" when X = 227 AND Y = 132 else
"000000000000" when X = 228 AND Y = 132 else
"000000000000" when X = 229 AND Y = 132 else
"000000000000" when X = 230 AND Y = 132 else
"000000000000" when X = 231 AND Y = 132 else
"000000000000" when X = 232 AND Y = 132 else
"000000000000" when X = 233 AND Y = 132 else
"000000000000" when X = 234 AND Y = 132 else
"000000000000" when X = 235 AND Y = 132 else
"000000000000" when X = 236 AND Y = 132 else
"000000000000" when X = 237 AND Y = 132 else
"000000000000" when X = 238 AND Y = 132 else
"000000000000" when X = 239 AND Y = 132 else
"000000000000" when X = 240 AND Y = 132 else
"000000000000" when X = 241 AND Y = 132 else
"000000000000" when X = 242 AND Y = 132 else
"000000000000" when X = 243 AND Y = 132 else
"000000000000" when X = 244 AND Y = 132 else
"000000000000" when X = 245 AND Y = 132 else
"000000000000" when X = 246 AND Y = 132 else
"000000000000" when X = 247 AND Y = 132 else
"000000000000" when X = 248 AND Y = 132 else
"000000000000" when X = 249 AND Y = 132 else
"000000000000" when X = 250 AND Y = 132 else
"000000000000" when X = 251 AND Y = 132 else
"000000000000" when X = 252 AND Y = 132 else
"000000000000" when X = 253 AND Y = 132 else
"000000000000" when X = 254 AND Y = 132 else
"000000000000" when X = 255 AND Y = 132 else
"000000000000" when X = 256 AND Y = 132 else
"000000000000" when X = 257 AND Y = 132 else
"000000000000" when X = 258 AND Y = 132 else
"000000000000" when X = 259 AND Y = 132 else
"000000000000" when X = 260 AND Y = 132 else
"000000000000" when X = 261 AND Y = 132 else
"000000000000" when X = 262 AND Y = 132 else
"000000000000" when X = 263 AND Y = 132 else
"000000000000" when X = 264 AND Y = 132 else
"000000000000" when X = 265 AND Y = 132 else
"000000000000" when X = 266 AND Y = 132 else
"000000000000" when X = 267 AND Y = 132 else
"000000000000" when X = 268 AND Y = 132 else
"000000000000" when X = 269 AND Y = 132 else
"000000000000" when X = 270 AND Y = 132 else
"000000000000" when X = 271 AND Y = 132 else
"000000000000" when X = 272 AND Y = 132 else
"000000000000" when X = 273 AND Y = 132 else
"000000000000" when X = 274 AND Y = 132 else
"000000000000" when X = 275 AND Y = 132 else
"000000000000" when X = 276 AND Y = 132 else
"000000000000" when X = 277 AND Y = 132 else
"000000000000" when X = 278 AND Y = 132 else
"000000000000" when X = 279 AND Y = 132 else
"000000000000" when X = 280 AND Y = 132 else
"000000000000" when X = 281 AND Y = 132 else
"000000000000" when X = 282 AND Y = 132 else
"000000000000" when X = 283 AND Y = 132 else
"000000000000" when X = 284 AND Y = 132 else
"000000000000" when X = 285 AND Y = 132 else
"000000000000" when X = 286 AND Y = 132 else
"000000000000" when X = 287 AND Y = 132 else
"000000000000" when X = 288 AND Y = 132 else
"000000000000" when X = 289 AND Y = 132 else
"000000000000" when X = 290 AND Y = 132 else
"000000000000" when X = 291 AND Y = 132 else
"000000000000" when X = 292 AND Y = 132 else
"000000000000" when X = 293 AND Y = 132 else
"000000000000" when X = 294 AND Y = 132 else
"000000000000" when X = 295 AND Y = 132 else
"000000000000" when X = 296 AND Y = 132 else
"000000000000" when X = 297 AND Y = 132 else
"000000000000" when X = 298 AND Y = 132 else
"000000000000" when X = 299 AND Y = 132 else
"000000000000" when X = 300 AND Y = 132 else
"000000000000" when X = 301 AND Y = 132 else
"000000000000" when X = 302 AND Y = 132 else
"000000000000" when X = 303 AND Y = 132 else
"000000000000" when X = 304 AND Y = 132 else
"000000000000" when X = 305 AND Y = 132 else
"000000000000" when X = 306 AND Y = 132 else
"000000000000" when X = 307 AND Y = 132 else
"000000000000" when X = 308 AND Y = 132 else
"000000000000" when X = 309 AND Y = 132 else
"000000000000" when X = 310 AND Y = 132 else
"000000000000" when X = 311 AND Y = 132 else
"000000000000" when X = 312 AND Y = 132 else
"000000000000" when X = 313 AND Y = 132 else
"000000000000" when X = 314 AND Y = 132 else
"000000000000" when X = 315 AND Y = 132 else
"000000000000" when X = 316 AND Y = 132 else
"000000000000" when X = 317 AND Y = 132 else
"000000000000" when X = 318 AND Y = 132 else
"000000000000" when X = 319 AND Y = 132 else
"000000000000" when X = 320 AND Y = 132 else
"000000000000" when X = 321 AND Y = 132 else
"000000000000" when X = 322 AND Y = 132 else
"000000000000" when X = 323 AND Y = 132 else
"000000000000" when X = 324 AND Y = 132 else
"000000000000" when X = 0 AND Y = 133 else
"000000000000" when X = 1 AND Y = 133 else
"000000000000" when X = 2 AND Y = 133 else
"000000000000" when X = 3 AND Y = 133 else
"000000000000" when X = 4 AND Y = 133 else
"000000000000" when X = 5 AND Y = 133 else
"000000000000" when X = 6 AND Y = 133 else
"000000000000" when X = 7 AND Y = 133 else
"000000000000" when X = 8 AND Y = 133 else
"000000000000" when X = 9 AND Y = 133 else
"000000000000" when X = 10 AND Y = 133 else
"000000000000" when X = 11 AND Y = 133 else
"000000000000" when X = 12 AND Y = 133 else
"000000000000" when X = 13 AND Y = 133 else
"000000000000" when X = 14 AND Y = 133 else
"000000000000" when X = 15 AND Y = 133 else
"000000000000" when X = 16 AND Y = 133 else
"000000000000" when X = 17 AND Y = 133 else
"000000000000" when X = 18 AND Y = 133 else
"000000000000" when X = 19 AND Y = 133 else
"000000000000" when X = 20 AND Y = 133 else
"000000000000" when X = 21 AND Y = 133 else
"000000000000" when X = 22 AND Y = 133 else
"000000000000" when X = 23 AND Y = 133 else
"000000000000" when X = 24 AND Y = 133 else
"000000000000" when X = 25 AND Y = 133 else
"000000000000" when X = 26 AND Y = 133 else
"000000000000" when X = 27 AND Y = 133 else
"000000000000" when X = 28 AND Y = 133 else
"000000000000" when X = 29 AND Y = 133 else
"000000000000" when X = 30 AND Y = 133 else
"000000000000" when X = 31 AND Y = 133 else
"000000000000" when X = 32 AND Y = 133 else
"000000000000" when X = 33 AND Y = 133 else
"000000000000" when X = 34 AND Y = 133 else
"000000000000" when X = 35 AND Y = 133 else
"000000000000" when X = 36 AND Y = 133 else
"000000000000" when X = 37 AND Y = 133 else
"000000000000" when X = 38 AND Y = 133 else
"000000000000" when X = 39 AND Y = 133 else
"100010011101" when X = 40 AND Y = 133 else
"100010011101" when X = 41 AND Y = 133 else
"100010011101" when X = 42 AND Y = 133 else
"100010011101" when X = 43 AND Y = 133 else
"100010011101" when X = 44 AND Y = 133 else
"100010011101" when X = 45 AND Y = 133 else
"100010011101" when X = 46 AND Y = 133 else
"100010011101" when X = 47 AND Y = 133 else
"100010011101" when X = 48 AND Y = 133 else
"100010011101" when X = 49 AND Y = 133 else
"100010011101" when X = 50 AND Y = 133 else
"100010011101" when X = 51 AND Y = 133 else
"100010011101" when X = 52 AND Y = 133 else
"100010011101" when X = 53 AND Y = 133 else
"100010011101" when X = 54 AND Y = 133 else
"100010011101" when X = 55 AND Y = 133 else
"100010011101" when X = 56 AND Y = 133 else
"100010011101" when X = 57 AND Y = 133 else
"100010011101" when X = 58 AND Y = 133 else
"100010011101" when X = 59 AND Y = 133 else
"100010011101" when X = 60 AND Y = 133 else
"100010011101" when X = 61 AND Y = 133 else
"100010011101" when X = 62 AND Y = 133 else
"100010011101" when X = 63 AND Y = 133 else
"100010011101" when X = 64 AND Y = 133 else
"100010011101" when X = 65 AND Y = 133 else
"100010011101" when X = 66 AND Y = 133 else
"100010011101" when X = 67 AND Y = 133 else
"100010011101" when X = 68 AND Y = 133 else
"100010011101" when X = 69 AND Y = 133 else
"100010011101" when X = 70 AND Y = 133 else
"100010011101" when X = 71 AND Y = 133 else
"100010011101" when X = 72 AND Y = 133 else
"100010011101" when X = 73 AND Y = 133 else
"100010011101" when X = 74 AND Y = 133 else
"100010011101" when X = 75 AND Y = 133 else
"100010011101" when X = 76 AND Y = 133 else
"100010011101" when X = 77 AND Y = 133 else
"100010011101" when X = 78 AND Y = 133 else
"100010011101" when X = 79 AND Y = 133 else
"100010011101" when X = 80 AND Y = 133 else
"100010011101" when X = 81 AND Y = 133 else
"100010011101" when X = 82 AND Y = 133 else
"100010011101" when X = 83 AND Y = 133 else
"100010011101" when X = 84 AND Y = 133 else
"100010011101" when X = 85 AND Y = 133 else
"100010011101" when X = 86 AND Y = 133 else
"100010011101" when X = 87 AND Y = 133 else
"100010011101" when X = 88 AND Y = 133 else
"100010011101" when X = 89 AND Y = 133 else
"100010011101" when X = 90 AND Y = 133 else
"100010011101" when X = 91 AND Y = 133 else
"100010011101" when X = 92 AND Y = 133 else
"100010011101" when X = 93 AND Y = 133 else
"100010011101" when X = 94 AND Y = 133 else
"100010011101" when X = 95 AND Y = 133 else
"100010011101" when X = 96 AND Y = 133 else
"100010011101" when X = 97 AND Y = 133 else
"100010011101" when X = 98 AND Y = 133 else
"100010011101" when X = 99 AND Y = 133 else
"100010011101" when X = 100 AND Y = 133 else
"100010011101" when X = 101 AND Y = 133 else
"100010011101" when X = 102 AND Y = 133 else
"100010011101" when X = 103 AND Y = 133 else
"100010011101" when X = 104 AND Y = 133 else
"100010011101" when X = 105 AND Y = 133 else
"100010011101" when X = 106 AND Y = 133 else
"100010011101" when X = 107 AND Y = 133 else
"100010011101" when X = 108 AND Y = 133 else
"100010011101" when X = 109 AND Y = 133 else
"110111011111" when X = 110 AND Y = 133 else
"110111011111" when X = 111 AND Y = 133 else
"110111011111" when X = 112 AND Y = 133 else
"110111011111" when X = 113 AND Y = 133 else
"110111011111" when X = 114 AND Y = 133 else
"110111011111" when X = 115 AND Y = 133 else
"110111011111" when X = 116 AND Y = 133 else
"110111011111" when X = 117 AND Y = 133 else
"110111011111" when X = 118 AND Y = 133 else
"110111011111" when X = 119 AND Y = 133 else
"110111011111" when X = 120 AND Y = 133 else
"110111011111" when X = 121 AND Y = 133 else
"110111011111" when X = 122 AND Y = 133 else
"110111011111" when X = 123 AND Y = 133 else
"110111011111" when X = 124 AND Y = 133 else
"110111011111" when X = 125 AND Y = 133 else
"110111011111" when X = 126 AND Y = 133 else
"110111011111" when X = 127 AND Y = 133 else
"110111011111" when X = 128 AND Y = 133 else
"110111011111" when X = 129 AND Y = 133 else
"110111011111" when X = 130 AND Y = 133 else
"110111011111" when X = 131 AND Y = 133 else
"110111011111" when X = 132 AND Y = 133 else
"110111011111" when X = 133 AND Y = 133 else
"110111011111" when X = 134 AND Y = 133 else
"110111011111" when X = 135 AND Y = 133 else
"110111011111" when X = 136 AND Y = 133 else
"110111011111" when X = 137 AND Y = 133 else
"110111011111" when X = 138 AND Y = 133 else
"110111011111" when X = 139 AND Y = 133 else
"110111011111" when X = 140 AND Y = 133 else
"110111011111" when X = 141 AND Y = 133 else
"110111011111" when X = 142 AND Y = 133 else
"110111011111" when X = 143 AND Y = 133 else
"110111011111" when X = 144 AND Y = 133 else
"110111011111" when X = 145 AND Y = 133 else
"110111011111" when X = 146 AND Y = 133 else
"110111011111" when X = 147 AND Y = 133 else
"110111011111" when X = 148 AND Y = 133 else
"110111011111" when X = 149 AND Y = 133 else
"110111011111" when X = 150 AND Y = 133 else
"110111011111" when X = 151 AND Y = 133 else
"110111011111" when X = 152 AND Y = 133 else
"110111011111" when X = 153 AND Y = 133 else
"110111011111" when X = 154 AND Y = 133 else
"110111011111" when X = 155 AND Y = 133 else
"110111011111" when X = 156 AND Y = 133 else
"110111011111" when X = 157 AND Y = 133 else
"110111011111" when X = 158 AND Y = 133 else
"110111011111" when X = 159 AND Y = 133 else
"110111011111" when X = 160 AND Y = 133 else
"110111011111" when X = 161 AND Y = 133 else
"110111011111" when X = 162 AND Y = 133 else
"110111011111" when X = 163 AND Y = 133 else
"110111011111" when X = 164 AND Y = 133 else
"110111011111" when X = 165 AND Y = 133 else
"110111011111" when X = 166 AND Y = 133 else
"110111011111" when X = 167 AND Y = 133 else
"110111011111" when X = 168 AND Y = 133 else
"110111011111" when X = 169 AND Y = 133 else
"110111011111" when X = 170 AND Y = 133 else
"110111011111" when X = 171 AND Y = 133 else
"110111011111" when X = 172 AND Y = 133 else
"110111011111" when X = 173 AND Y = 133 else
"110111011111" when X = 174 AND Y = 133 else
"110111011111" when X = 175 AND Y = 133 else
"110111011111" when X = 176 AND Y = 133 else
"110111011111" when X = 177 AND Y = 133 else
"110111011111" when X = 178 AND Y = 133 else
"110111011111" when X = 179 AND Y = 133 else
"110111011111" when X = 180 AND Y = 133 else
"110111011111" when X = 181 AND Y = 133 else
"110111011111" when X = 182 AND Y = 133 else
"110111011111" when X = 183 AND Y = 133 else
"110111011111" when X = 184 AND Y = 133 else
"110111011111" when X = 185 AND Y = 133 else
"110111011111" when X = 186 AND Y = 133 else
"110111011111" when X = 187 AND Y = 133 else
"110111011111" when X = 188 AND Y = 133 else
"110111011111" when X = 189 AND Y = 133 else
"110111011111" when X = 190 AND Y = 133 else
"110111011111" when X = 191 AND Y = 133 else
"110111011111" when X = 192 AND Y = 133 else
"110111011111" when X = 193 AND Y = 133 else
"110111011111" when X = 194 AND Y = 133 else
"110111011111" when X = 195 AND Y = 133 else
"110111011111" when X = 196 AND Y = 133 else
"110111011111" when X = 197 AND Y = 133 else
"110111011111" when X = 198 AND Y = 133 else
"110111011111" when X = 199 AND Y = 133 else
"000000000000" when X = 200 AND Y = 133 else
"000000000000" when X = 201 AND Y = 133 else
"000000000000" when X = 202 AND Y = 133 else
"000000000000" when X = 203 AND Y = 133 else
"000000000000" when X = 204 AND Y = 133 else
"000000000000" when X = 205 AND Y = 133 else
"000000000000" when X = 206 AND Y = 133 else
"000000000000" when X = 207 AND Y = 133 else
"000000000000" when X = 208 AND Y = 133 else
"000000000000" when X = 209 AND Y = 133 else
"000000000000" when X = 210 AND Y = 133 else
"000000000000" when X = 211 AND Y = 133 else
"000000000000" when X = 212 AND Y = 133 else
"000000000000" when X = 213 AND Y = 133 else
"000000000000" when X = 214 AND Y = 133 else
"000000000000" when X = 215 AND Y = 133 else
"000000000000" when X = 216 AND Y = 133 else
"000000000000" when X = 217 AND Y = 133 else
"000000000000" when X = 218 AND Y = 133 else
"000000000000" when X = 219 AND Y = 133 else
"000000000000" when X = 220 AND Y = 133 else
"000000000000" when X = 221 AND Y = 133 else
"000000000000" when X = 222 AND Y = 133 else
"000000000000" when X = 223 AND Y = 133 else
"000000000000" when X = 224 AND Y = 133 else
"000000000000" when X = 225 AND Y = 133 else
"000000000000" when X = 226 AND Y = 133 else
"000000000000" when X = 227 AND Y = 133 else
"000000000000" when X = 228 AND Y = 133 else
"000000000000" when X = 229 AND Y = 133 else
"000000000000" when X = 230 AND Y = 133 else
"000000000000" when X = 231 AND Y = 133 else
"000000000000" when X = 232 AND Y = 133 else
"000000000000" when X = 233 AND Y = 133 else
"000000000000" when X = 234 AND Y = 133 else
"000000000000" when X = 235 AND Y = 133 else
"000000000000" when X = 236 AND Y = 133 else
"000000000000" when X = 237 AND Y = 133 else
"000000000000" when X = 238 AND Y = 133 else
"000000000000" when X = 239 AND Y = 133 else
"000000000000" when X = 240 AND Y = 133 else
"000000000000" when X = 241 AND Y = 133 else
"000000000000" when X = 242 AND Y = 133 else
"000000000000" when X = 243 AND Y = 133 else
"000000000000" when X = 244 AND Y = 133 else
"000000000000" when X = 245 AND Y = 133 else
"000000000000" when X = 246 AND Y = 133 else
"000000000000" when X = 247 AND Y = 133 else
"000000000000" when X = 248 AND Y = 133 else
"000000000000" when X = 249 AND Y = 133 else
"000000000000" when X = 250 AND Y = 133 else
"000000000000" when X = 251 AND Y = 133 else
"000000000000" when X = 252 AND Y = 133 else
"000000000000" when X = 253 AND Y = 133 else
"000000000000" when X = 254 AND Y = 133 else
"000000000000" when X = 255 AND Y = 133 else
"000000000000" when X = 256 AND Y = 133 else
"000000000000" when X = 257 AND Y = 133 else
"000000000000" when X = 258 AND Y = 133 else
"000000000000" when X = 259 AND Y = 133 else
"000000000000" when X = 260 AND Y = 133 else
"000000000000" when X = 261 AND Y = 133 else
"000000000000" when X = 262 AND Y = 133 else
"000000000000" when X = 263 AND Y = 133 else
"000000000000" when X = 264 AND Y = 133 else
"000000000000" when X = 265 AND Y = 133 else
"000000000000" when X = 266 AND Y = 133 else
"000000000000" when X = 267 AND Y = 133 else
"000000000000" when X = 268 AND Y = 133 else
"000000000000" when X = 269 AND Y = 133 else
"000000000000" when X = 270 AND Y = 133 else
"000000000000" when X = 271 AND Y = 133 else
"000000000000" when X = 272 AND Y = 133 else
"000000000000" when X = 273 AND Y = 133 else
"000000000000" when X = 274 AND Y = 133 else
"000000000000" when X = 275 AND Y = 133 else
"000000000000" when X = 276 AND Y = 133 else
"000000000000" when X = 277 AND Y = 133 else
"000000000000" when X = 278 AND Y = 133 else
"000000000000" when X = 279 AND Y = 133 else
"000000000000" when X = 280 AND Y = 133 else
"000000000000" when X = 281 AND Y = 133 else
"000000000000" when X = 282 AND Y = 133 else
"000000000000" when X = 283 AND Y = 133 else
"000000000000" when X = 284 AND Y = 133 else
"000000000000" when X = 285 AND Y = 133 else
"000000000000" when X = 286 AND Y = 133 else
"000000000000" when X = 287 AND Y = 133 else
"000000000000" when X = 288 AND Y = 133 else
"000000000000" when X = 289 AND Y = 133 else
"000000000000" when X = 290 AND Y = 133 else
"000000000000" when X = 291 AND Y = 133 else
"000000000000" when X = 292 AND Y = 133 else
"000000000000" when X = 293 AND Y = 133 else
"000000000000" when X = 294 AND Y = 133 else
"000000000000" when X = 295 AND Y = 133 else
"000000000000" when X = 296 AND Y = 133 else
"000000000000" when X = 297 AND Y = 133 else
"000000000000" when X = 298 AND Y = 133 else
"000000000000" when X = 299 AND Y = 133 else
"000000000000" when X = 300 AND Y = 133 else
"000000000000" when X = 301 AND Y = 133 else
"000000000000" when X = 302 AND Y = 133 else
"000000000000" when X = 303 AND Y = 133 else
"000000000000" when X = 304 AND Y = 133 else
"000000000000" when X = 305 AND Y = 133 else
"000000000000" when X = 306 AND Y = 133 else
"000000000000" when X = 307 AND Y = 133 else
"000000000000" when X = 308 AND Y = 133 else
"000000000000" when X = 309 AND Y = 133 else
"000000000000" when X = 310 AND Y = 133 else
"000000000000" when X = 311 AND Y = 133 else
"000000000000" when X = 312 AND Y = 133 else
"000000000000" when X = 313 AND Y = 133 else
"000000000000" when X = 314 AND Y = 133 else
"000000000000" when X = 315 AND Y = 133 else
"000000000000" when X = 316 AND Y = 133 else
"000000000000" when X = 317 AND Y = 133 else
"000000000000" when X = 318 AND Y = 133 else
"000000000000" when X = 319 AND Y = 133 else
"000000000000" when X = 320 AND Y = 133 else
"000000000000" when X = 321 AND Y = 133 else
"000000000000" when X = 322 AND Y = 133 else
"000000000000" when X = 323 AND Y = 133 else
"000000000000" when X = 324 AND Y = 133 else
"000000000000" when X = 0 AND Y = 134 else
"000000000000" when X = 1 AND Y = 134 else
"000000000000" when X = 2 AND Y = 134 else
"000000000000" when X = 3 AND Y = 134 else
"000000000000" when X = 4 AND Y = 134 else
"000000000000" when X = 5 AND Y = 134 else
"000000000000" when X = 6 AND Y = 134 else
"000000000000" when X = 7 AND Y = 134 else
"000000000000" when X = 8 AND Y = 134 else
"000000000000" when X = 9 AND Y = 134 else
"000000000000" when X = 10 AND Y = 134 else
"000000000000" when X = 11 AND Y = 134 else
"000000000000" when X = 12 AND Y = 134 else
"000000000000" when X = 13 AND Y = 134 else
"000000000000" when X = 14 AND Y = 134 else
"000000000000" when X = 15 AND Y = 134 else
"000000000000" when X = 16 AND Y = 134 else
"000000000000" when X = 17 AND Y = 134 else
"000000000000" when X = 18 AND Y = 134 else
"000000000000" when X = 19 AND Y = 134 else
"000000000000" when X = 20 AND Y = 134 else
"000000000000" when X = 21 AND Y = 134 else
"000000000000" when X = 22 AND Y = 134 else
"000000000000" when X = 23 AND Y = 134 else
"000000000000" when X = 24 AND Y = 134 else
"000000000000" when X = 25 AND Y = 134 else
"000000000000" when X = 26 AND Y = 134 else
"000000000000" when X = 27 AND Y = 134 else
"000000000000" when X = 28 AND Y = 134 else
"000000000000" when X = 29 AND Y = 134 else
"000000000000" when X = 30 AND Y = 134 else
"000000000000" when X = 31 AND Y = 134 else
"000000000000" when X = 32 AND Y = 134 else
"000000000000" when X = 33 AND Y = 134 else
"000000000000" when X = 34 AND Y = 134 else
"000000000000" when X = 35 AND Y = 134 else
"000000000000" when X = 36 AND Y = 134 else
"000000000000" when X = 37 AND Y = 134 else
"000000000000" when X = 38 AND Y = 134 else
"000000000000" when X = 39 AND Y = 134 else
"100010011101" when X = 40 AND Y = 134 else
"100010011101" when X = 41 AND Y = 134 else
"100010011101" when X = 42 AND Y = 134 else
"100010011101" when X = 43 AND Y = 134 else
"100010011101" when X = 44 AND Y = 134 else
"100010011101" when X = 45 AND Y = 134 else
"100010011101" when X = 46 AND Y = 134 else
"100010011101" when X = 47 AND Y = 134 else
"100010011101" when X = 48 AND Y = 134 else
"100010011101" when X = 49 AND Y = 134 else
"100010011101" when X = 50 AND Y = 134 else
"100010011101" when X = 51 AND Y = 134 else
"100010011101" when X = 52 AND Y = 134 else
"100010011101" when X = 53 AND Y = 134 else
"100010011101" when X = 54 AND Y = 134 else
"100010011101" when X = 55 AND Y = 134 else
"100010011101" when X = 56 AND Y = 134 else
"100010011101" when X = 57 AND Y = 134 else
"100010011101" when X = 58 AND Y = 134 else
"100010011101" when X = 59 AND Y = 134 else
"100010011101" when X = 60 AND Y = 134 else
"100010011101" when X = 61 AND Y = 134 else
"100010011101" when X = 62 AND Y = 134 else
"100010011101" when X = 63 AND Y = 134 else
"100010011101" when X = 64 AND Y = 134 else
"100010011101" when X = 65 AND Y = 134 else
"100010011101" when X = 66 AND Y = 134 else
"100010011101" when X = 67 AND Y = 134 else
"100010011101" when X = 68 AND Y = 134 else
"100010011101" when X = 69 AND Y = 134 else
"100010011101" when X = 70 AND Y = 134 else
"100010011101" when X = 71 AND Y = 134 else
"100010011101" when X = 72 AND Y = 134 else
"100010011101" when X = 73 AND Y = 134 else
"100010011101" when X = 74 AND Y = 134 else
"100010011101" when X = 75 AND Y = 134 else
"100010011101" when X = 76 AND Y = 134 else
"100010011101" when X = 77 AND Y = 134 else
"100010011101" when X = 78 AND Y = 134 else
"100010011101" when X = 79 AND Y = 134 else
"100010011101" when X = 80 AND Y = 134 else
"100010011101" when X = 81 AND Y = 134 else
"100010011101" when X = 82 AND Y = 134 else
"100010011101" when X = 83 AND Y = 134 else
"100010011101" when X = 84 AND Y = 134 else
"100010011101" when X = 85 AND Y = 134 else
"100010011101" when X = 86 AND Y = 134 else
"100010011101" when X = 87 AND Y = 134 else
"100010011101" when X = 88 AND Y = 134 else
"100010011101" when X = 89 AND Y = 134 else
"100010011101" when X = 90 AND Y = 134 else
"100010011101" when X = 91 AND Y = 134 else
"100010011101" when X = 92 AND Y = 134 else
"100010011101" when X = 93 AND Y = 134 else
"100010011101" when X = 94 AND Y = 134 else
"100010011101" when X = 95 AND Y = 134 else
"100010011101" when X = 96 AND Y = 134 else
"100010011101" when X = 97 AND Y = 134 else
"100010011101" when X = 98 AND Y = 134 else
"100010011101" when X = 99 AND Y = 134 else
"100010011101" when X = 100 AND Y = 134 else
"100010011101" when X = 101 AND Y = 134 else
"100010011101" when X = 102 AND Y = 134 else
"100010011101" when X = 103 AND Y = 134 else
"100010011101" when X = 104 AND Y = 134 else
"100010011101" when X = 105 AND Y = 134 else
"100010011101" when X = 106 AND Y = 134 else
"100010011101" when X = 107 AND Y = 134 else
"100010011101" when X = 108 AND Y = 134 else
"100010011101" when X = 109 AND Y = 134 else
"110111011111" when X = 110 AND Y = 134 else
"110111011111" when X = 111 AND Y = 134 else
"110111011111" when X = 112 AND Y = 134 else
"110111011111" when X = 113 AND Y = 134 else
"110111011111" when X = 114 AND Y = 134 else
"110111011111" when X = 115 AND Y = 134 else
"110111011111" when X = 116 AND Y = 134 else
"110111011111" when X = 117 AND Y = 134 else
"110111011111" when X = 118 AND Y = 134 else
"110111011111" when X = 119 AND Y = 134 else
"110111011111" when X = 120 AND Y = 134 else
"110111011111" when X = 121 AND Y = 134 else
"110111011111" when X = 122 AND Y = 134 else
"110111011111" when X = 123 AND Y = 134 else
"110111011111" when X = 124 AND Y = 134 else
"110111011111" when X = 125 AND Y = 134 else
"110111011111" when X = 126 AND Y = 134 else
"110111011111" when X = 127 AND Y = 134 else
"110111011111" when X = 128 AND Y = 134 else
"110111011111" when X = 129 AND Y = 134 else
"110111011111" when X = 130 AND Y = 134 else
"110111011111" when X = 131 AND Y = 134 else
"110111011111" when X = 132 AND Y = 134 else
"110111011111" when X = 133 AND Y = 134 else
"110111011111" when X = 134 AND Y = 134 else
"110111011111" when X = 135 AND Y = 134 else
"110111011111" when X = 136 AND Y = 134 else
"110111011111" when X = 137 AND Y = 134 else
"110111011111" when X = 138 AND Y = 134 else
"110111011111" when X = 139 AND Y = 134 else
"110111011111" when X = 140 AND Y = 134 else
"110111011111" when X = 141 AND Y = 134 else
"110111011111" when X = 142 AND Y = 134 else
"110111011111" when X = 143 AND Y = 134 else
"110111011111" when X = 144 AND Y = 134 else
"110111011111" when X = 145 AND Y = 134 else
"110111011111" when X = 146 AND Y = 134 else
"110111011111" when X = 147 AND Y = 134 else
"110111011111" when X = 148 AND Y = 134 else
"110111011111" when X = 149 AND Y = 134 else
"110111011111" when X = 150 AND Y = 134 else
"110111011111" when X = 151 AND Y = 134 else
"110111011111" when X = 152 AND Y = 134 else
"110111011111" when X = 153 AND Y = 134 else
"110111011111" when X = 154 AND Y = 134 else
"110111011111" when X = 155 AND Y = 134 else
"110111011111" when X = 156 AND Y = 134 else
"110111011111" when X = 157 AND Y = 134 else
"110111011111" when X = 158 AND Y = 134 else
"110111011111" when X = 159 AND Y = 134 else
"110111011111" when X = 160 AND Y = 134 else
"110111011111" when X = 161 AND Y = 134 else
"110111011111" when X = 162 AND Y = 134 else
"110111011111" when X = 163 AND Y = 134 else
"110111011111" when X = 164 AND Y = 134 else
"110111011111" when X = 165 AND Y = 134 else
"110111011111" when X = 166 AND Y = 134 else
"110111011111" when X = 167 AND Y = 134 else
"110111011111" when X = 168 AND Y = 134 else
"110111011111" when X = 169 AND Y = 134 else
"110111011111" when X = 170 AND Y = 134 else
"110111011111" when X = 171 AND Y = 134 else
"110111011111" when X = 172 AND Y = 134 else
"110111011111" when X = 173 AND Y = 134 else
"110111011111" when X = 174 AND Y = 134 else
"110111011111" when X = 175 AND Y = 134 else
"110111011111" when X = 176 AND Y = 134 else
"110111011111" when X = 177 AND Y = 134 else
"110111011111" when X = 178 AND Y = 134 else
"110111011111" when X = 179 AND Y = 134 else
"110111011111" when X = 180 AND Y = 134 else
"110111011111" when X = 181 AND Y = 134 else
"110111011111" when X = 182 AND Y = 134 else
"110111011111" when X = 183 AND Y = 134 else
"110111011111" when X = 184 AND Y = 134 else
"110111011111" when X = 185 AND Y = 134 else
"110111011111" when X = 186 AND Y = 134 else
"110111011111" when X = 187 AND Y = 134 else
"110111011111" when X = 188 AND Y = 134 else
"110111011111" when X = 189 AND Y = 134 else
"110111011111" when X = 190 AND Y = 134 else
"110111011111" when X = 191 AND Y = 134 else
"110111011111" when X = 192 AND Y = 134 else
"110111011111" when X = 193 AND Y = 134 else
"110111011111" when X = 194 AND Y = 134 else
"110111011111" when X = 195 AND Y = 134 else
"110111011111" when X = 196 AND Y = 134 else
"110111011111" when X = 197 AND Y = 134 else
"110111011111" when X = 198 AND Y = 134 else
"110111011111" when X = 199 AND Y = 134 else
"000000000000" when X = 200 AND Y = 134 else
"000000000000" when X = 201 AND Y = 134 else
"000000000000" when X = 202 AND Y = 134 else
"000000000000" when X = 203 AND Y = 134 else
"000000000000" when X = 204 AND Y = 134 else
"000000000000" when X = 205 AND Y = 134 else
"000000000000" when X = 206 AND Y = 134 else
"000000000000" when X = 207 AND Y = 134 else
"000000000000" when X = 208 AND Y = 134 else
"000000000000" when X = 209 AND Y = 134 else
"000000000000" when X = 210 AND Y = 134 else
"000000000000" when X = 211 AND Y = 134 else
"000000000000" when X = 212 AND Y = 134 else
"000000000000" when X = 213 AND Y = 134 else
"000000000000" when X = 214 AND Y = 134 else
"000000000000" when X = 215 AND Y = 134 else
"000000000000" when X = 216 AND Y = 134 else
"000000000000" when X = 217 AND Y = 134 else
"000000000000" when X = 218 AND Y = 134 else
"000000000000" when X = 219 AND Y = 134 else
"000000000000" when X = 220 AND Y = 134 else
"000000000000" when X = 221 AND Y = 134 else
"000000000000" when X = 222 AND Y = 134 else
"000000000000" when X = 223 AND Y = 134 else
"000000000000" when X = 224 AND Y = 134 else
"000000000000" when X = 225 AND Y = 134 else
"000000000000" when X = 226 AND Y = 134 else
"000000000000" when X = 227 AND Y = 134 else
"000000000000" when X = 228 AND Y = 134 else
"000000000000" when X = 229 AND Y = 134 else
"000000000000" when X = 230 AND Y = 134 else
"000000000000" when X = 231 AND Y = 134 else
"000000000000" when X = 232 AND Y = 134 else
"000000000000" when X = 233 AND Y = 134 else
"000000000000" when X = 234 AND Y = 134 else
"000000000000" when X = 235 AND Y = 134 else
"000000000000" when X = 236 AND Y = 134 else
"000000000000" when X = 237 AND Y = 134 else
"000000000000" when X = 238 AND Y = 134 else
"000000000000" when X = 239 AND Y = 134 else
"000000000000" when X = 240 AND Y = 134 else
"000000000000" when X = 241 AND Y = 134 else
"000000000000" when X = 242 AND Y = 134 else
"000000000000" when X = 243 AND Y = 134 else
"000000000000" when X = 244 AND Y = 134 else
"000000000000" when X = 245 AND Y = 134 else
"000000000000" when X = 246 AND Y = 134 else
"000000000000" when X = 247 AND Y = 134 else
"000000000000" when X = 248 AND Y = 134 else
"000000000000" when X = 249 AND Y = 134 else
"000000000000" when X = 250 AND Y = 134 else
"000000000000" when X = 251 AND Y = 134 else
"000000000000" when X = 252 AND Y = 134 else
"000000000000" when X = 253 AND Y = 134 else
"000000000000" when X = 254 AND Y = 134 else
"000000000000" when X = 255 AND Y = 134 else
"000000000000" when X = 256 AND Y = 134 else
"000000000000" when X = 257 AND Y = 134 else
"000000000000" when X = 258 AND Y = 134 else
"000000000000" when X = 259 AND Y = 134 else
"000000000000" when X = 260 AND Y = 134 else
"000000000000" when X = 261 AND Y = 134 else
"000000000000" when X = 262 AND Y = 134 else
"000000000000" when X = 263 AND Y = 134 else
"000000000000" when X = 264 AND Y = 134 else
"000000000000" when X = 265 AND Y = 134 else
"000000000000" when X = 266 AND Y = 134 else
"000000000000" when X = 267 AND Y = 134 else
"000000000000" when X = 268 AND Y = 134 else
"000000000000" when X = 269 AND Y = 134 else
"000000000000" when X = 270 AND Y = 134 else
"000000000000" when X = 271 AND Y = 134 else
"000000000000" when X = 272 AND Y = 134 else
"000000000000" when X = 273 AND Y = 134 else
"000000000000" when X = 274 AND Y = 134 else
"000000000000" when X = 275 AND Y = 134 else
"000000000000" when X = 276 AND Y = 134 else
"000000000000" when X = 277 AND Y = 134 else
"000000000000" when X = 278 AND Y = 134 else
"000000000000" when X = 279 AND Y = 134 else
"000000000000" when X = 280 AND Y = 134 else
"000000000000" when X = 281 AND Y = 134 else
"000000000000" when X = 282 AND Y = 134 else
"000000000000" when X = 283 AND Y = 134 else
"000000000000" when X = 284 AND Y = 134 else
"000000000000" when X = 285 AND Y = 134 else
"000000000000" when X = 286 AND Y = 134 else
"000000000000" when X = 287 AND Y = 134 else
"000000000000" when X = 288 AND Y = 134 else
"000000000000" when X = 289 AND Y = 134 else
"000000000000" when X = 290 AND Y = 134 else
"000000000000" when X = 291 AND Y = 134 else
"000000000000" when X = 292 AND Y = 134 else
"000000000000" when X = 293 AND Y = 134 else
"000000000000" when X = 294 AND Y = 134 else
"000000000000" when X = 295 AND Y = 134 else
"000000000000" when X = 296 AND Y = 134 else
"000000000000" when X = 297 AND Y = 134 else
"000000000000" when X = 298 AND Y = 134 else
"000000000000" when X = 299 AND Y = 134 else
"000000000000" when X = 300 AND Y = 134 else
"000000000000" when X = 301 AND Y = 134 else
"000000000000" when X = 302 AND Y = 134 else
"000000000000" when X = 303 AND Y = 134 else
"000000000000" when X = 304 AND Y = 134 else
"000000000000" when X = 305 AND Y = 134 else
"000000000000" when X = 306 AND Y = 134 else
"000000000000" when X = 307 AND Y = 134 else
"000000000000" when X = 308 AND Y = 134 else
"000000000000" when X = 309 AND Y = 134 else
"000000000000" when X = 310 AND Y = 134 else
"000000000000" when X = 311 AND Y = 134 else
"000000000000" when X = 312 AND Y = 134 else
"000000000000" when X = 313 AND Y = 134 else
"000000000000" when X = 314 AND Y = 134 else
"000000000000" when X = 315 AND Y = 134 else
"000000000000" when X = 316 AND Y = 134 else
"000000000000" when X = 317 AND Y = 134 else
"000000000000" when X = 318 AND Y = 134 else
"000000000000" when X = 319 AND Y = 134 else
"000000000000" when X = 320 AND Y = 134 else
"000000000000" when X = 321 AND Y = 134 else
"000000000000" when X = 322 AND Y = 134 else
"000000000000" when X = 323 AND Y = 134 else
"000000000000" when X = 324 AND Y = 134 else
"000000000000"; -- should never get here
end rtl;
