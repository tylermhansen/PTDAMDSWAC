-- Tyler Hansen
-- CS232 Final Project
-- genSpriteROM.py
-- generates a ROM file in VHDL from a .ppm image

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity road_texture is
port(
X	: in INTEGER RANGE 0 TO 1688;
Y	: in INTEGER RANGE 0 TO 1688;
data : out std_logic_vector (11 downto 0)
);

end entity;

architecture rtl of road_texture is
begin
data <=
"111000100000" when X = 0 AND Y = 0 else
"111000100000" when X = 1 AND Y = 0 else
"111000100000" when X = 2 AND Y = 0 else
"111000100000" when X = 3 AND Y = 0 else
"111000100000" when X = 4 AND Y = 0 else
"111000100000" when X = 5 AND Y = 0 else
"111000100000" when X = 6 AND Y = 0 else
"111000100000" when X = 7 AND Y = 0 else
"111000100000" when X = 8 AND Y = 0 else
"111000100000" when X = 9 AND Y = 0 else
"111000100000" when X = 10 AND Y = 0 else
"111000100000" when X = 11 AND Y = 0 else
"111000100000" when X = 12 AND Y = 0 else
"111000100000" when X = 13 AND Y = 0 else
"111000100000" when X = 14 AND Y = 0 else
"111000100000" when X = 15 AND Y = 0 else
"010101010101" when X = 16 AND Y = 0 else
"010101010101" when X = 17 AND Y = 0 else
"010101010101" when X = 18 AND Y = 0 else
"010101010101" when X = 19 AND Y = 0 else
"010101010101" when X = 20 AND Y = 0 else
"010101010101" when X = 21 AND Y = 0 else
"010101010101" when X = 22 AND Y = 0 else
"010101010101" when X = 23 AND Y = 0 else
"010101010101" when X = 24 AND Y = 0 else
"111011101110" when X = 25 AND Y = 0 else
"111011101110" when X = 26 AND Y = 0 else
"111011101110" when X = 27 AND Y = 0 else
"111011101110" when X = 28 AND Y = 0 else
"010101010101" when X = 29 AND Y = 0 else
"010101010101" when X = 30 AND Y = 0 else
"010101010101" when X = 31 AND Y = 0 else
"010101010101" when X = 32 AND Y = 0 else
"010101010101" when X = 33 AND Y = 0 else
"010101010101" when X = 34 AND Y = 0 else
"010101010101" when X = 35 AND Y = 0 else
"010101010101" when X = 36 AND Y = 0 else
"010101010101" when X = 37 AND Y = 0 else
"010101010101" when X = 38 AND Y = 0 else
"010101010101" when X = 39 AND Y = 0 else
"010101010101" when X = 40 AND Y = 0 else
"010101010101" when X = 41 AND Y = 0 else
"010101010101" when X = 42 AND Y = 0 else
"010101010101" when X = 43 AND Y = 0 else
"010101010101" when X = 44 AND Y = 0 else
"010101010101" when X = 45 AND Y = 0 else
"010101010101" when X = 46 AND Y = 0 else
"010101010101" when X = 47 AND Y = 0 else
"010101010101" when X = 48 AND Y = 0 else
"010101010101" when X = 49 AND Y = 0 else
"010101010101" when X = 50 AND Y = 0 else
"010101010101" when X = 51 AND Y = 0 else
"010101010101" when X = 52 AND Y = 0 else
"010101010101" when X = 53 AND Y = 0 else
"010101010101" when X = 54 AND Y = 0 else
"010101010101" when X = 55 AND Y = 0 else
"010101010101" when X = 56 AND Y = 0 else
"010101010101" when X = 57 AND Y = 0 else
"010101010101" when X = 58 AND Y = 0 else
"010101010101" when X = 59 AND Y = 0 else
"010101010101" when X = 60 AND Y = 0 else
"010101010101" when X = 61 AND Y = 0 else
"010101010101" when X = 62 AND Y = 0 else
"010101010101" when X = 63 AND Y = 0 else
"010101010101" when X = 64 AND Y = 0 else
"010101010101" when X = 65 AND Y = 0 else
"010101010101" when X = 66 AND Y = 0 else
"010101010101" when X = 67 AND Y = 0 else
"010101010101" when X = 68 AND Y = 0 else
"010101010101" when X = 69 AND Y = 0 else
"010101010101" when X = 70 AND Y = 0 else
"010101010101" when X = 71 AND Y = 0 else
"010101010101" when X = 72 AND Y = 0 else
"010101010101" when X = 73 AND Y = 0 else
"010101010101" when X = 74 AND Y = 0 else
"010101010101" when X = 75 AND Y = 0 else
"010101010101" when X = 76 AND Y = 0 else
"010101010101" when X = 77 AND Y = 0 else
"010101010101" when X = 78 AND Y = 0 else
"010101010101" when X = 79 AND Y = 0 else
"010101010101" when X = 80 AND Y = 0 else
"010101010101" when X = 81 AND Y = 0 else
"010101010101" when X = 82 AND Y = 0 else
"010101010101" when X = 83 AND Y = 0 else
"010101010101" when X = 84 AND Y = 0 else
"010101010101" when X = 85 AND Y = 0 else
"010101010101" when X = 86 AND Y = 0 else
"010101010101" when X = 87 AND Y = 0 else
"010101010101" when X = 88 AND Y = 0 else
"010101010101" when X = 89 AND Y = 0 else
"010101010101" when X = 90 AND Y = 0 else
"010101010101" when X = 91 AND Y = 0 else
"010101010101" when X = 92 AND Y = 0 else
"010101010101" when X = 93 AND Y = 0 else
"010101010101" when X = 94 AND Y = 0 else
"010101010101" when X = 95 AND Y = 0 else
"010101010101" when X = 96 AND Y = 0 else
"010101010101" when X = 97 AND Y = 0 else
"010101010101" when X = 98 AND Y = 0 else
"010101010101" when X = 99 AND Y = 0 else
"010101010101" when X = 100 AND Y = 0 else
"010101010101" when X = 101 AND Y = 0 else
"010101010101" when X = 102 AND Y = 0 else
"010101010101" when X = 103 AND Y = 0 else
"010101010101" when X = 104 AND Y = 0 else
"010101010101" when X = 105 AND Y = 0 else
"010101010101" when X = 106 AND Y = 0 else
"010101010101" when X = 107 AND Y = 0 else
"010101010101" when X = 108 AND Y = 0 else
"010101010101" when X = 109 AND Y = 0 else
"010101010101" when X = 110 AND Y = 0 else
"010101010101" when X = 111 AND Y = 0 else
"010101010101" when X = 112 AND Y = 0 else
"010101010101" when X = 113 AND Y = 0 else
"010101010101" when X = 114 AND Y = 0 else
"010101010101" when X = 115 AND Y = 0 else
"010101010101" when X = 116 AND Y = 0 else
"010101010101" when X = 117 AND Y = 0 else
"010101010101" when X = 118 AND Y = 0 else
"010101010101" when X = 119 AND Y = 0 else
"010101010101" when X = 120 AND Y = 0 else
"010101010101" when X = 121 AND Y = 0 else
"010101010101" when X = 122 AND Y = 0 else
"010101010101" when X = 123 AND Y = 0 else
"010101010101" when X = 124 AND Y = 0 else
"010101010101" when X = 125 AND Y = 0 else
"111011101110" when X = 126 AND Y = 0 else
"111011101110" when X = 127 AND Y = 0 else
"111011101110" when X = 128 AND Y = 0 else
"111011101110" when X = 129 AND Y = 0 else
"010101010101" when X = 130 AND Y = 0 else
"010101010101" when X = 131 AND Y = 0 else
"010101010101" when X = 132 AND Y = 0 else
"010101010101" when X = 133 AND Y = 0 else
"010101010101" when X = 134 AND Y = 0 else
"010101010101" when X = 135 AND Y = 0 else
"010101010101" when X = 136 AND Y = 0 else
"010101010101" when X = 137 AND Y = 0 else
"010101010101" when X = 138 AND Y = 0 else
"010101010101" when X = 139 AND Y = 0 else
"010101010101" when X = 140 AND Y = 0 else
"010101010101" when X = 141 AND Y = 0 else
"010101010101" when X = 142 AND Y = 0 else
"010101010101" when X = 143 AND Y = 0 else
"010101010101" when X = 144 AND Y = 0 else
"010101010101" when X = 145 AND Y = 0 else
"010101010101" when X = 146 AND Y = 0 else
"010101010101" when X = 147 AND Y = 0 else
"010101010101" when X = 148 AND Y = 0 else
"010101010101" when X = 149 AND Y = 0 else
"010101010101" when X = 150 AND Y = 0 else
"010101010101" when X = 151 AND Y = 0 else
"010101010101" when X = 152 AND Y = 0 else
"010101010101" when X = 153 AND Y = 0 else
"010101010101" when X = 154 AND Y = 0 else
"010101010101" when X = 155 AND Y = 0 else
"010101010101" when X = 156 AND Y = 0 else
"010101010101" when X = 157 AND Y = 0 else
"010101010101" when X = 158 AND Y = 0 else
"010101010101" when X = 159 AND Y = 0 else
"010101010101" when X = 160 AND Y = 0 else
"010101010101" when X = 161 AND Y = 0 else
"010101010101" when X = 162 AND Y = 0 else
"010101010101" when X = 163 AND Y = 0 else
"010101010101" when X = 164 AND Y = 0 else
"010101010101" when X = 165 AND Y = 0 else
"010101010101" when X = 166 AND Y = 0 else
"010101010101" when X = 167 AND Y = 0 else
"010101010101" when X = 168 AND Y = 0 else
"010101010101" when X = 169 AND Y = 0 else
"010101010101" when X = 170 AND Y = 0 else
"010101010101" when X = 171 AND Y = 0 else
"010101010101" when X = 172 AND Y = 0 else
"010101010101" when X = 173 AND Y = 0 else
"010101010101" when X = 174 AND Y = 0 else
"010101010101" when X = 175 AND Y = 0 else
"010101010101" when X = 176 AND Y = 0 else
"010101010101" when X = 177 AND Y = 0 else
"010101010101" when X = 178 AND Y = 0 else
"010101010101" when X = 179 AND Y = 0 else
"010101010101" when X = 180 AND Y = 0 else
"010101010101" when X = 181 AND Y = 0 else
"010101010101" when X = 182 AND Y = 0 else
"010101010101" when X = 183 AND Y = 0 else
"010101010101" when X = 184 AND Y = 0 else
"010101010101" when X = 185 AND Y = 0 else
"010101010101" when X = 186 AND Y = 0 else
"010101010101" when X = 187 AND Y = 0 else
"010101010101" when X = 188 AND Y = 0 else
"010101010101" when X = 189 AND Y = 0 else
"010101010101" when X = 190 AND Y = 0 else
"010101010101" when X = 191 AND Y = 0 else
"010101010101" when X = 192 AND Y = 0 else
"010101010101" when X = 193 AND Y = 0 else
"010101010101" when X = 194 AND Y = 0 else
"010101010101" when X = 195 AND Y = 0 else
"010101010101" when X = 196 AND Y = 0 else
"010101010101" when X = 197 AND Y = 0 else
"010101010101" when X = 198 AND Y = 0 else
"010101010101" when X = 199 AND Y = 0 else
"010101010101" when X = 200 AND Y = 0 else
"010101010101" when X = 201 AND Y = 0 else
"010101010101" when X = 202 AND Y = 0 else
"010101010101" when X = 203 AND Y = 0 else
"010101010101" when X = 204 AND Y = 0 else
"010101010101" when X = 205 AND Y = 0 else
"010101010101" when X = 206 AND Y = 0 else
"010101010101" when X = 207 AND Y = 0 else
"010101010101" when X = 208 AND Y = 0 else
"010101010101" when X = 209 AND Y = 0 else
"010101010101" when X = 210 AND Y = 0 else
"010101010101" when X = 211 AND Y = 0 else
"010101010101" when X = 212 AND Y = 0 else
"010101010101" when X = 213 AND Y = 0 else
"010101010101" when X = 214 AND Y = 0 else
"010101010101" when X = 215 AND Y = 0 else
"010101010101" when X = 216 AND Y = 0 else
"010101010101" when X = 217 AND Y = 0 else
"010101010101" when X = 218 AND Y = 0 else
"010101010101" when X = 219 AND Y = 0 else
"010101010101" when X = 220 AND Y = 0 else
"010101010101" when X = 221 AND Y = 0 else
"010101010101" when X = 222 AND Y = 0 else
"010101010101" when X = 223 AND Y = 0 else
"010101010101" when X = 224 AND Y = 0 else
"010101010101" when X = 225 AND Y = 0 else
"010101010101" when X = 226 AND Y = 0 else
"111011101110" when X = 227 AND Y = 0 else
"111011101110" when X = 228 AND Y = 0 else
"111011101110" when X = 229 AND Y = 0 else
"111011101110" when X = 230 AND Y = 0 else
"010101010101" when X = 231 AND Y = 0 else
"010101010101" when X = 232 AND Y = 0 else
"010101010101" when X = 233 AND Y = 0 else
"010101010101" when X = 234 AND Y = 0 else
"010101010101" when X = 235 AND Y = 0 else
"010101010101" when X = 236 AND Y = 0 else
"010101010101" when X = 237 AND Y = 0 else
"010101010101" when X = 238 AND Y = 0 else
"010101010101" when X = 239 AND Y = 0 else
"111000100000" when X = 240 AND Y = 0 else
"111000100000" when X = 241 AND Y = 0 else
"111000100000" when X = 242 AND Y = 0 else
"111000100000" when X = 243 AND Y = 0 else
"111000100000" when X = 244 AND Y = 0 else
"111000100000" when X = 245 AND Y = 0 else
"111000100000" when X = 246 AND Y = 0 else
"111000100000" when X = 247 AND Y = 0 else
"111000100000" when X = 248 AND Y = 0 else
"111000100000" when X = 249 AND Y = 0 else
"111000100000" when X = 250 AND Y = 0 else
"111000100000" when X = 251 AND Y = 0 else
"111000100000" when X = 252 AND Y = 0 else
"111000100000" when X = 253 AND Y = 0 else
"111000100000" when X = 254 AND Y = 0 else
"111000100000" when X = 255 AND Y = 0 else
"111011101110" when X = 0 AND Y = 1 else
"111011101110" when X = 1 AND Y = 1 else
"111011101110" when X = 2 AND Y = 1 else
"111011101110" when X = 3 AND Y = 1 else
"111011101110" when X = 4 AND Y = 1 else
"111011101110" when X = 5 AND Y = 1 else
"111011101110" when X = 6 AND Y = 1 else
"111011101110" when X = 7 AND Y = 1 else
"111011101110" when X = 8 AND Y = 1 else
"111011101110" when X = 9 AND Y = 1 else
"111011101110" when X = 10 AND Y = 1 else
"111011101110" when X = 11 AND Y = 1 else
"111011101110" when X = 12 AND Y = 1 else
"111011101110" when X = 13 AND Y = 1 else
"111011101110" when X = 14 AND Y = 1 else
"111011101110" when X = 15 AND Y = 1 else
"010101010101" when X = 16 AND Y = 1 else
"010101010101" when X = 17 AND Y = 1 else
"010101010101" when X = 18 AND Y = 1 else
"010101010101" when X = 19 AND Y = 1 else
"010101010101" when X = 20 AND Y = 1 else
"010101010101" when X = 21 AND Y = 1 else
"010101010101" when X = 22 AND Y = 1 else
"010101010101" when X = 23 AND Y = 1 else
"010101010101" when X = 24 AND Y = 1 else
"111011101110" when X = 25 AND Y = 1 else
"111011101110" when X = 26 AND Y = 1 else
"111011101110" when X = 27 AND Y = 1 else
"111011101110" when X = 28 AND Y = 1 else
"010101010101" when X = 29 AND Y = 1 else
"010101010101" when X = 30 AND Y = 1 else
"010101010101" when X = 31 AND Y = 1 else
"010101010101" when X = 32 AND Y = 1 else
"010101010101" when X = 33 AND Y = 1 else
"010101010101" when X = 34 AND Y = 1 else
"010101010101" when X = 35 AND Y = 1 else
"010101010101" when X = 36 AND Y = 1 else
"010101010101" when X = 37 AND Y = 1 else
"010101010101" when X = 38 AND Y = 1 else
"010101010101" when X = 39 AND Y = 1 else
"010101010101" when X = 40 AND Y = 1 else
"010101010101" when X = 41 AND Y = 1 else
"010101010101" when X = 42 AND Y = 1 else
"010101010101" when X = 43 AND Y = 1 else
"010101010101" when X = 44 AND Y = 1 else
"010101010101" when X = 45 AND Y = 1 else
"010101010101" when X = 46 AND Y = 1 else
"010101010101" when X = 47 AND Y = 1 else
"010101010101" when X = 48 AND Y = 1 else
"010101010101" when X = 49 AND Y = 1 else
"010101010101" when X = 50 AND Y = 1 else
"010101010101" when X = 51 AND Y = 1 else
"010101010101" when X = 52 AND Y = 1 else
"010101010101" when X = 53 AND Y = 1 else
"010101010101" when X = 54 AND Y = 1 else
"010101010101" when X = 55 AND Y = 1 else
"010101010101" when X = 56 AND Y = 1 else
"010101010101" when X = 57 AND Y = 1 else
"010101010101" when X = 58 AND Y = 1 else
"010101010101" when X = 59 AND Y = 1 else
"010101010101" when X = 60 AND Y = 1 else
"010101010101" when X = 61 AND Y = 1 else
"010101010101" when X = 62 AND Y = 1 else
"010101010101" when X = 63 AND Y = 1 else
"010101010101" when X = 64 AND Y = 1 else
"010101010101" when X = 65 AND Y = 1 else
"010101010101" when X = 66 AND Y = 1 else
"010101010101" when X = 67 AND Y = 1 else
"010101010101" when X = 68 AND Y = 1 else
"010101010101" when X = 69 AND Y = 1 else
"010101010101" when X = 70 AND Y = 1 else
"010101010101" when X = 71 AND Y = 1 else
"010101010101" when X = 72 AND Y = 1 else
"010101010101" when X = 73 AND Y = 1 else
"010101010101" when X = 74 AND Y = 1 else
"010101010101" when X = 75 AND Y = 1 else
"010101010101" when X = 76 AND Y = 1 else
"010101010101" when X = 77 AND Y = 1 else
"010101010101" when X = 78 AND Y = 1 else
"010101010101" when X = 79 AND Y = 1 else
"010101010101" when X = 80 AND Y = 1 else
"010101010101" when X = 81 AND Y = 1 else
"010101010101" when X = 82 AND Y = 1 else
"010101010101" when X = 83 AND Y = 1 else
"010101010101" when X = 84 AND Y = 1 else
"010101010101" when X = 85 AND Y = 1 else
"010101010101" when X = 86 AND Y = 1 else
"010101010101" when X = 87 AND Y = 1 else
"010101010101" when X = 88 AND Y = 1 else
"010101010101" when X = 89 AND Y = 1 else
"010101010101" when X = 90 AND Y = 1 else
"010101010101" when X = 91 AND Y = 1 else
"010101010101" when X = 92 AND Y = 1 else
"010101010101" when X = 93 AND Y = 1 else
"010101010101" when X = 94 AND Y = 1 else
"010101010101" when X = 95 AND Y = 1 else
"010101010101" when X = 96 AND Y = 1 else
"010101010101" when X = 97 AND Y = 1 else
"010101010101" when X = 98 AND Y = 1 else
"010101010101" when X = 99 AND Y = 1 else
"010101010101" when X = 100 AND Y = 1 else
"010101010101" when X = 101 AND Y = 1 else
"010101010101" when X = 102 AND Y = 1 else
"010101010101" when X = 103 AND Y = 1 else
"010101010101" when X = 104 AND Y = 1 else
"010101010101" when X = 105 AND Y = 1 else
"010101010101" when X = 106 AND Y = 1 else
"010101010101" when X = 107 AND Y = 1 else
"010101010101" when X = 108 AND Y = 1 else
"010101010101" when X = 109 AND Y = 1 else
"010101010101" when X = 110 AND Y = 1 else
"010101010101" when X = 111 AND Y = 1 else
"010101010101" when X = 112 AND Y = 1 else
"010101010101" when X = 113 AND Y = 1 else
"010101010101" when X = 114 AND Y = 1 else
"010101010101" when X = 115 AND Y = 1 else
"010101010101" when X = 116 AND Y = 1 else
"010101010101" when X = 117 AND Y = 1 else
"010101010101" when X = 118 AND Y = 1 else
"010101010101" when X = 119 AND Y = 1 else
"010101010101" when X = 120 AND Y = 1 else
"010101010101" when X = 121 AND Y = 1 else
"010101010101" when X = 122 AND Y = 1 else
"010101010101" when X = 123 AND Y = 1 else
"010101010101" when X = 124 AND Y = 1 else
"010101010101" when X = 125 AND Y = 1 else
"111011101110" when X = 126 AND Y = 1 else
"111011101110" when X = 127 AND Y = 1 else
"111011101110" when X = 128 AND Y = 1 else
"111011101110" when X = 129 AND Y = 1 else
"010101010101" when X = 130 AND Y = 1 else
"010101010101" when X = 131 AND Y = 1 else
"010101010101" when X = 132 AND Y = 1 else
"010101010101" when X = 133 AND Y = 1 else
"010101010101" when X = 134 AND Y = 1 else
"010101010101" when X = 135 AND Y = 1 else
"010101010101" when X = 136 AND Y = 1 else
"010101010101" when X = 137 AND Y = 1 else
"010101010101" when X = 138 AND Y = 1 else
"010101010101" when X = 139 AND Y = 1 else
"010101010101" when X = 140 AND Y = 1 else
"010101010101" when X = 141 AND Y = 1 else
"010101010101" when X = 142 AND Y = 1 else
"010101010101" when X = 143 AND Y = 1 else
"010101010101" when X = 144 AND Y = 1 else
"010101010101" when X = 145 AND Y = 1 else
"010101010101" when X = 146 AND Y = 1 else
"010101010101" when X = 147 AND Y = 1 else
"010101010101" when X = 148 AND Y = 1 else
"010101010101" when X = 149 AND Y = 1 else
"010101010101" when X = 150 AND Y = 1 else
"010101010101" when X = 151 AND Y = 1 else
"010101010101" when X = 152 AND Y = 1 else
"010101010101" when X = 153 AND Y = 1 else
"010101010101" when X = 154 AND Y = 1 else
"010101010101" when X = 155 AND Y = 1 else
"010101010101" when X = 156 AND Y = 1 else
"010101010101" when X = 157 AND Y = 1 else
"010101010101" when X = 158 AND Y = 1 else
"010101010101" when X = 159 AND Y = 1 else
"010101010101" when X = 160 AND Y = 1 else
"010101010101" when X = 161 AND Y = 1 else
"010101010101" when X = 162 AND Y = 1 else
"010101010101" when X = 163 AND Y = 1 else
"010101010101" when X = 164 AND Y = 1 else
"010101010101" when X = 165 AND Y = 1 else
"010101010101" when X = 166 AND Y = 1 else
"010101010101" when X = 167 AND Y = 1 else
"010101010101" when X = 168 AND Y = 1 else
"010101010101" when X = 169 AND Y = 1 else
"010101010101" when X = 170 AND Y = 1 else
"010101010101" when X = 171 AND Y = 1 else
"010101010101" when X = 172 AND Y = 1 else
"010101010101" when X = 173 AND Y = 1 else
"010101010101" when X = 174 AND Y = 1 else
"010101010101" when X = 175 AND Y = 1 else
"010101010101" when X = 176 AND Y = 1 else
"010101010101" when X = 177 AND Y = 1 else
"010101010101" when X = 178 AND Y = 1 else
"010101010101" when X = 179 AND Y = 1 else
"010101010101" when X = 180 AND Y = 1 else
"010101010101" when X = 181 AND Y = 1 else
"010101010101" when X = 182 AND Y = 1 else
"010101010101" when X = 183 AND Y = 1 else
"010101010101" when X = 184 AND Y = 1 else
"010101010101" when X = 185 AND Y = 1 else
"010101010101" when X = 186 AND Y = 1 else
"010101010101" when X = 187 AND Y = 1 else
"010101010101" when X = 188 AND Y = 1 else
"010101010101" when X = 189 AND Y = 1 else
"010101010101" when X = 190 AND Y = 1 else
"010101010101" when X = 191 AND Y = 1 else
"010101010101" when X = 192 AND Y = 1 else
"010101010101" when X = 193 AND Y = 1 else
"010101010101" when X = 194 AND Y = 1 else
"010101010101" when X = 195 AND Y = 1 else
"010101010101" when X = 196 AND Y = 1 else
"010101010101" when X = 197 AND Y = 1 else
"010101010101" when X = 198 AND Y = 1 else
"010101010101" when X = 199 AND Y = 1 else
"010101010101" when X = 200 AND Y = 1 else
"010101010101" when X = 201 AND Y = 1 else
"010101010101" when X = 202 AND Y = 1 else
"010101010101" when X = 203 AND Y = 1 else
"010101010101" when X = 204 AND Y = 1 else
"010101010101" when X = 205 AND Y = 1 else
"010101010101" when X = 206 AND Y = 1 else
"010101010101" when X = 207 AND Y = 1 else
"010101010101" when X = 208 AND Y = 1 else
"010101010101" when X = 209 AND Y = 1 else
"010101010101" when X = 210 AND Y = 1 else
"010101010101" when X = 211 AND Y = 1 else
"010101010101" when X = 212 AND Y = 1 else
"010101010101" when X = 213 AND Y = 1 else
"010101010101" when X = 214 AND Y = 1 else
"010101010101" when X = 215 AND Y = 1 else
"010101010101" when X = 216 AND Y = 1 else
"010101010101" when X = 217 AND Y = 1 else
"010101010101" when X = 218 AND Y = 1 else
"010101010101" when X = 219 AND Y = 1 else
"010101010101" when X = 220 AND Y = 1 else
"010101010101" when X = 221 AND Y = 1 else
"010101010101" when X = 222 AND Y = 1 else
"010101010101" when X = 223 AND Y = 1 else
"010101010101" when X = 224 AND Y = 1 else
"010101010101" when X = 225 AND Y = 1 else
"010101010101" when X = 226 AND Y = 1 else
"111011101110" when X = 227 AND Y = 1 else
"111011101110" when X = 228 AND Y = 1 else
"111011101110" when X = 229 AND Y = 1 else
"111011101110" when X = 230 AND Y = 1 else
"010101010101" when X = 231 AND Y = 1 else
"010101010101" when X = 232 AND Y = 1 else
"010101010101" when X = 233 AND Y = 1 else
"010101010101" when X = 234 AND Y = 1 else
"010101010101" when X = 235 AND Y = 1 else
"010101010101" when X = 236 AND Y = 1 else
"010101010101" when X = 237 AND Y = 1 else
"010101010101" when X = 238 AND Y = 1 else
"010101010101" when X = 239 AND Y = 1 else
"111011101110" when X = 240 AND Y = 1 else
"111011101110" when X = 241 AND Y = 1 else
"111011101110" when X = 242 AND Y = 1 else
"111011101110" when X = 243 AND Y = 1 else
"111011101110" when X = 244 AND Y = 1 else
"111011101110" when X = 245 AND Y = 1 else
"111011101110" when X = 246 AND Y = 1 else
"111011101110" when X = 247 AND Y = 1 else
"111011101110" when X = 248 AND Y = 1 else
"111011101110" when X = 249 AND Y = 1 else
"111011101110" when X = 250 AND Y = 1 else
"111011101110" when X = 251 AND Y = 1 else
"111011101110" when X = 252 AND Y = 1 else
"111011101110" when X = 253 AND Y = 1 else
"111011101110" when X = 254 AND Y = 1 else
"111011101110" when X = 255 AND Y = 1 else
"111000100000" when X = 0 AND Y = 2 else
"111000100000" when X = 1 AND Y = 2 else
"111000100000" when X = 2 AND Y = 2 else
"111000100000" when X = 3 AND Y = 2 else
"111000100000" when X = 4 AND Y = 2 else
"111000100000" when X = 5 AND Y = 2 else
"111000100000" when X = 6 AND Y = 2 else
"111000100000" when X = 7 AND Y = 2 else
"111000100000" when X = 8 AND Y = 2 else
"111000100000" when X = 9 AND Y = 2 else
"111000100000" when X = 10 AND Y = 2 else
"111000100000" when X = 11 AND Y = 2 else
"111000100000" when X = 12 AND Y = 2 else
"111000100000" when X = 13 AND Y = 2 else
"111000100000" when X = 14 AND Y = 2 else
"111000100000" when X = 15 AND Y = 2 else
"010101010101" when X = 16 AND Y = 2 else
"010101010101" when X = 17 AND Y = 2 else
"010101010101" when X = 18 AND Y = 2 else
"010101010101" when X = 19 AND Y = 2 else
"010101010101" when X = 20 AND Y = 2 else
"010101010101" when X = 21 AND Y = 2 else
"010101010101" when X = 22 AND Y = 2 else
"010101010101" when X = 23 AND Y = 2 else
"010101010101" when X = 24 AND Y = 2 else
"111011101110" when X = 25 AND Y = 2 else
"111011101110" when X = 26 AND Y = 2 else
"111011101110" when X = 27 AND Y = 2 else
"111011101110" when X = 28 AND Y = 2 else
"010101010101" when X = 29 AND Y = 2 else
"010101010101" when X = 30 AND Y = 2 else
"010101010101" when X = 31 AND Y = 2 else
"010101010101" when X = 32 AND Y = 2 else
"010101010101" when X = 33 AND Y = 2 else
"010101010101" when X = 34 AND Y = 2 else
"010101010101" when X = 35 AND Y = 2 else
"010101010101" when X = 36 AND Y = 2 else
"010101010101" when X = 37 AND Y = 2 else
"010101010101" when X = 38 AND Y = 2 else
"010101010101" when X = 39 AND Y = 2 else
"010101010101" when X = 40 AND Y = 2 else
"010101010101" when X = 41 AND Y = 2 else
"010101010101" when X = 42 AND Y = 2 else
"010101010101" when X = 43 AND Y = 2 else
"010101010101" when X = 44 AND Y = 2 else
"010101010101" when X = 45 AND Y = 2 else
"010101010101" when X = 46 AND Y = 2 else
"010101010101" when X = 47 AND Y = 2 else
"010101010101" when X = 48 AND Y = 2 else
"010101010101" when X = 49 AND Y = 2 else
"010101010101" when X = 50 AND Y = 2 else
"010101010101" when X = 51 AND Y = 2 else
"010101010101" when X = 52 AND Y = 2 else
"010101010101" when X = 53 AND Y = 2 else
"010101010101" when X = 54 AND Y = 2 else
"010101010101" when X = 55 AND Y = 2 else
"010101010101" when X = 56 AND Y = 2 else
"010101010101" when X = 57 AND Y = 2 else
"010101010101" when X = 58 AND Y = 2 else
"010101010101" when X = 59 AND Y = 2 else
"010101010101" when X = 60 AND Y = 2 else
"010101010101" when X = 61 AND Y = 2 else
"010101010101" when X = 62 AND Y = 2 else
"010101010101" when X = 63 AND Y = 2 else
"010101010101" when X = 64 AND Y = 2 else
"010101010101" when X = 65 AND Y = 2 else
"010101010101" when X = 66 AND Y = 2 else
"010101010101" when X = 67 AND Y = 2 else
"010101010101" when X = 68 AND Y = 2 else
"010101010101" when X = 69 AND Y = 2 else
"010101010101" when X = 70 AND Y = 2 else
"010101010101" when X = 71 AND Y = 2 else
"010101010101" when X = 72 AND Y = 2 else
"010101010101" when X = 73 AND Y = 2 else
"010101010101" when X = 74 AND Y = 2 else
"010101010101" when X = 75 AND Y = 2 else
"010101010101" when X = 76 AND Y = 2 else
"010101010101" when X = 77 AND Y = 2 else
"010101010101" when X = 78 AND Y = 2 else
"010101010101" when X = 79 AND Y = 2 else
"010101010101" when X = 80 AND Y = 2 else
"010101010101" when X = 81 AND Y = 2 else
"010101010101" when X = 82 AND Y = 2 else
"010101010101" when X = 83 AND Y = 2 else
"010101010101" when X = 84 AND Y = 2 else
"010101010101" when X = 85 AND Y = 2 else
"010101010101" when X = 86 AND Y = 2 else
"010101010101" when X = 87 AND Y = 2 else
"010101010101" when X = 88 AND Y = 2 else
"010101010101" when X = 89 AND Y = 2 else
"010101010101" when X = 90 AND Y = 2 else
"010101010101" when X = 91 AND Y = 2 else
"010101010101" when X = 92 AND Y = 2 else
"010101010101" when X = 93 AND Y = 2 else
"010101010101" when X = 94 AND Y = 2 else
"010101010101" when X = 95 AND Y = 2 else
"010101010101" when X = 96 AND Y = 2 else
"010101010101" when X = 97 AND Y = 2 else
"010101010101" when X = 98 AND Y = 2 else
"010101010101" when X = 99 AND Y = 2 else
"010101010101" when X = 100 AND Y = 2 else
"010101010101" when X = 101 AND Y = 2 else
"010101010101" when X = 102 AND Y = 2 else
"010101010101" when X = 103 AND Y = 2 else
"010101010101" when X = 104 AND Y = 2 else
"010101010101" when X = 105 AND Y = 2 else
"010101010101" when X = 106 AND Y = 2 else
"010101010101" when X = 107 AND Y = 2 else
"010101010101" when X = 108 AND Y = 2 else
"010101010101" when X = 109 AND Y = 2 else
"010101010101" when X = 110 AND Y = 2 else
"010101010101" when X = 111 AND Y = 2 else
"010101010101" when X = 112 AND Y = 2 else
"010101010101" when X = 113 AND Y = 2 else
"010101010101" when X = 114 AND Y = 2 else
"010101010101" when X = 115 AND Y = 2 else
"010101010101" when X = 116 AND Y = 2 else
"010101010101" when X = 117 AND Y = 2 else
"010101010101" when X = 118 AND Y = 2 else
"010101010101" when X = 119 AND Y = 2 else
"010101010101" when X = 120 AND Y = 2 else
"010101010101" when X = 121 AND Y = 2 else
"010101010101" when X = 122 AND Y = 2 else
"010101010101" when X = 123 AND Y = 2 else
"010101010101" when X = 124 AND Y = 2 else
"010101010101" when X = 125 AND Y = 2 else
"010101010101" when X = 126 AND Y = 2 else
"010101010101" when X = 127 AND Y = 2 else
"010101010101" when X = 128 AND Y = 2 else
"010101010101" when X = 129 AND Y = 2 else
"010101010101" when X = 130 AND Y = 2 else
"010101010101" when X = 131 AND Y = 2 else
"010101010101" when X = 132 AND Y = 2 else
"010101010101" when X = 133 AND Y = 2 else
"010101010101" when X = 134 AND Y = 2 else
"010101010101" when X = 135 AND Y = 2 else
"010101010101" when X = 136 AND Y = 2 else
"010101010101" when X = 137 AND Y = 2 else
"010101010101" when X = 138 AND Y = 2 else
"010101010101" when X = 139 AND Y = 2 else
"010101010101" when X = 140 AND Y = 2 else
"010101010101" when X = 141 AND Y = 2 else
"010101010101" when X = 142 AND Y = 2 else
"010101010101" when X = 143 AND Y = 2 else
"010101010101" when X = 144 AND Y = 2 else
"010101010101" when X = 145 AND Y = 2 else
"010101010101" when X = 146 AND Y = 2 else
"010101010101" when X = 147 AND Y = 2 else
"010101010101" when X = 148 AND Y = 2 else
"010101010101" when X = 149 AND Y = 2 else
"010101010101" when X = 150 AND Y = 2 else
"010101010101" when X = 151 AND Y = 2 else
"010101010101" when X = 152 AND Y = 2 else
"010101010101" when X = 153 AND Y = 2 else
"010101010101" when X = 154 AND Y = 2 else
"010101010101" when X = 155 AND Y = 2 else
"010101010101" when X = 156 AND Y = 2 else
"010101010101" when X = 157 AND Y = 2 else
"010101010101" when X = 158 AND Y = 2 else
"010101010101" when X = 159 AND Y = 2 else
"010101010101" when X = 160 AND Y = 2 else
"010101010101" when X = 161 AND Y = 2 else
"010101010101" when X = 162 AND Y = 2 else
"010101010101" when X = 163 AND Y = 2 else
"010101010101" when X = 164 AND Y = 2 else
"010101010101" when X = 165 AND Y = 2 else
"010101010101" when X = 166 AND Y = 2 else
"010101010101" when X = 167 AND Y = 2 else
"010101010101" when X = 168 AND Y = 2 else
"010101010101" when X = 169 AND Y = 2 else
"010101010101" when X = 170 AND Y = 2 else
"010101010101" when X = 171 AND Y = 2 else
"010101010101" when X = 172 AND Y = 2 else
"010101010101" when X = 173 AND Y = 2 else
"010101010101" when X = 174 AND Y = 2 else
"010101010101" when X = 175 AND Y = 2 else
"010101010101" when X = 176 AND Y = 2 else
"010101010101" when X = 177 AND Y = 2 else
"010101010101" when X = 178 AND Y = 2 else
"010101010101" when X = 179 AND Y = 2 else
"010101010101" when X = 180 AND Y = 2 else
"010101010101" when X = 181 AND Y = 2 else
"010101010101" when X = 182 AND Y = 2 else
"010101010101" when X = 183 AND Y = 2 else
"010101010101" when X = 184 AND Y = 2 else
"010101010101" when X = 185 AND Y = 2 else
"010101010101" when X = 186 AND Y = 2 else
"010101010101" when X = 187 AND Y = 2 else
"010101010101" when X = 188 AND Y = 2 else
"010101010101" when X = 189 AND Y = 2 else
"010101010101" when X = 190 AND Y = 2 else
"010101010101" when X = 191 AND Y = 2 else
"010101010101" when X = 192 AND Y = 2 else
"010101010101" when X = 193 AND Y = 2 else
"010101010101" when X = 194 AND Y = 2 else
"010101010101" when X = 195 AND Y = 2 else
"010101010101" when X = 196 AND Y = 2 else
"010101010101" when X = 197 AND Y = 2 else
"010101010101" when X = 198 AND Y = 2 else
"010101010101" when X = 199 AND Y = 2 else
"010101010101" when X = 200 AND Y = 2 else
"010101010101" when X = 201 AND Y = 2 else
"010101010101" when X = 202 AND Y = 2 else
"010101010101" when X = 203 AND Y = 2 else
"010101010101" when X = 204 AND Y = 2 else
"010101010101" when X = 205 AND Y = 2 else
"010101010101" when X = 206 AND Y = 2 else
"010101010101" when X = 207 AND Y = 2 else
"010101010101" when X = 208 AND Y = 2 else
"010101010101" when X = 209 AND Y = 2 else
"010101010101" when X = 210 AND Y = 2 else
"010101010101" when X = 211 AND Y = 2 else
"010101010101" when X = 212 AND Y = 2 else
"010101010101" when X = 213 AND Y = 2 else
"010101010101" when X = 214 AND Y = 2 else
"010101010101" when X = 215 AND Y = 2 else
"010101010101" when X = 216 AND Y = 2 else
"010101010101" when X = 217 AND Y = 2 else
"010101010101" when X = 218 AND Y = 2 else
"010101010101" when X = 219 AND Y = 2 else
"010101010101" when X = 220 AND Y = 2 else
"010101010101" when X = 221 AND Y = 2 else
"010101010101" when X = 222 AND Y = 2 else
"010101010101" when X = 223 AND Y = 2 else
"010101010101" when X = 224 AND Y = 2 else
"010101010101" when X = 225 AND Y = 2 else
"010101010101" when X = 226 AND Y = 2 else
"111011101110" when X = 227 AND Y = 2 else
"111011101110" when X = 228 AND Y = 2 else
"111011101110" when X = 229 AND Y = 2 else
"111011101110" when X = 230 AND Y = 2 else
"010101010101" when X = 231 AND Y = 2 else
"010101010101" when X = 232 AND Y = 2 else
"010101010101" when X = 233 AND Y = 2 else
"010101010101" when X = 234 AND Y = 2 else
"010101010101" when X = 235 AND Y = 2 else
"010101010101" when X = 236 AND Y = 2 else
"010101010101" when X = 237 AND Y = 2 else
"010101010101" when X = 238 AND Y = 2 else
"010101010101" when X = 239 AND Y = 2 else
"111000100000" when X = 240 AND Y = 2 else
"111000100000" when X = 241 AND Y = 2 else
"111000100000" when X = 242 AND Y = 2 else
"111000100000" when X = 243 AND Y = 2 else
"111000100000" when X = 244 AND Y = 2 else
"111000100000" when X = 245 AND Y = 2 else
"111000100000" when X = 246 AND Y = 2 else
"111000100000" when X = 247 AND Y = 2 else
"111000100000" when X = 248 AND Y = 2 else
"111000100000" when X = 249 AND Y = 2 else
"111000100000" when X = 250 AND Y = 2 else
"111000100000" when X = 251 AND Y = 2 else
"111000100000" when X = 252 AND Y = 2 else
"111000100000" when X = 253 AND Y = 2 else
"111000100000" when X = 254 AND Y = 2 else
"111000100000" when X = 255 AND Y = 2 else
"111011101110" when X = 0 AND Y = 3 else
"111011101110" when X = 1 AND Y = 3 else
"111011101110" when X = 2 AND Y = 3 else
"111011101110" when X = 3 AND Y = 3 else
"111011101110" when X = 4 AND Y = 3 else
"111011101110" when X = 5 AND Y = 3 else
"111011101110" when X = 6 AND Y = 3 else
"111011101110" when X = 7 AND Y = 3 else
"111011101110" when X = 8 AND Y = 3 else
"111011101110" when X = 9 AND Y = 3 else
"111011101110" when X = 10 AND Y = 3 else
"111011101110" when X = 11 AND Y = 3 else
"111011101110" when X = 12 AND Y = 3 else
"111011101110" when X = 13 AND Y = 3 else
"111011101110" when X = 14 AND Y = 3 else
"111011101110" when X = 15 AND Y = 3 else
"010101010101" when X = 16 AND Y = 3 else
"010101010101" when X = 17 AND Y = 3 else
"010101010101" when X = 18 AND Y = 3 else
"010101010101" when X = 19 AND Y = 3 else
"010101010101" when X = 20 AND Y = 3 else
"010101010101" when X = 21 AND Y = 3 else
"010101010101" when X = 22 AND Y = 3 else
"010101010101" when X = 23 AND Y = 3 else
"010101010101" when X = 24 AND Y = 3 else
"111011101110" when X = 25 AND Y = 3 else
"111011101110" when X = 26 AND Y = 3 else
"111011101110" when X = 27 AND Y = 3 else
"111011101110" when X = 28 AND Y = 3 else
"010101010101" when X = 29 AND Y = 3 else
"010101010101" when X = 30 AND Y = 3 else
"010101010101" when X = 31 AND Y = 3 else
"010101010101" when X = 32 AND Y = 3 else
"010101010101" when X = 33 AND Y = 3 else
"010101010101" when X = 34 AND Y = 3 else
"010101010101" when X = 35 AND Y = 3 else
"010101010101" when X = 36 AND Y = 3 else
"010101010101" when X = 37 AND Y = 3 else
"010101010101" when X = 38 AND Y = 3 else
"010101010101" when X = 39 AND Y = 3 else
"010101010101" when X = 40 AND Y = 3 else
"010101010101" when X = 41 AND Y = 3 else
"010101010101" when X = 42 AND Y = 3 else
"010101010101" when X = 43 AND Y = 3 else
"010101010101" when X = 44 AND Y = 3 else
"010101010101" when X = 45 AND Y = 3 else
"010101010101" when X = 46 AND Y = 3 else
"010101010101" when X = 47 AND Y = 3 else
"010101010101" when X = 48 AND Y = 3 else
"010101010101" when X = 49 AND Y = 3 else
"010101010101" when X = 50 AND Y = 3 else
"010101010101" when X = 51 AND Y = 3 else
"010101010101" when X = 52 AND Y = 3 else
"010101010101" when X = 53 AND Y = 3 else
"010101010101" when X = 54 AND Y = 3 else
"010101010101" when X = 55 AND Y = 3 else
"010101010101" when X = 56 AND Y = 3 else
"010101010101" when X = 57 AND Y = 3 else
"010101010101" when X = 58 AND Y = 3 else
"010101010101" when X = 59 AND Y = 3 else
"010101010101" when X = 60 AND Y = 3 else
"010101010101" when X = 61 AND Y = 3 else
"010101010101" when X = 62 AND Y = 3 else
"010101010101" when X = 63 AND Y = 3 else
"010101010101" when X = 64 AND Y = 3 else
"010101010101" when X = 65 AND Y = 3 else
"010101010101" when X = 66 AND Y = 3 else
"010101010101" when X = 67 AND Y = 3 else
"010101010101" when X = 68 AND Y = 3 else
"010101010101" when X = 69 AND Y = 3 else
"010101010101" when X = 70 AND Y = 3 else
"010101010101" when X = 71 AND Y = 3 else
"010101010101" when X = 72 AND Y = 3 else
"010101010101" when X = 73 AND Y = 3 else
"010101010101" when X = 74 AND Y = 3 else
"010101010101" when X = 75 AND Y = 3 else
"010101010101" when X = 76 AND Y = 3 else
"010101010101" when X = 77 AND Y = 3 else
"010101010101" when X = 78 AND Y = 3 else
"010101010101" when X = 79 AND Y = 3 else
"010101010101" when X = 80 AND Y = 3 else
"010101010101" when X = 81 AND Y = 3 else
"010101010101" when X = 82 AND Y = 3 else
"010101010101" when X = 83 AND Y = 3 else
"010101010101" when X = 84 AND Y = 3 else
"010101010101" when X = 85 AND Y = 3 else
"010101010101" when X = 86 AND Y = 3 else
"010101010101" when X = 87 AND Y = 3 else
"010101010101" when X = 88 AND Y = 3 else
"010101010101" when X = 89 AND Y = 3 else
"010101010101" when X = 90 AND Y = 3 else
"010101010101" when X = 91 AND Y = 3 else
"010101010101" when X = 92 AND Y = 3 else
"010101010101" when X = 93 AND Y = 3 else
"010101010101" when X = 94 AND Y = 3 else
"010101010101" when X = 95 AND Y = 3 else
"010101010101" when X = 96 AND Y = 3 else
"010101010101" when X = 97 AND Y = 3 else
"010101010101" when X = 98 AND Y = 3 else
"010101010101" when X = 99 AND Y = 3 else
"010101010101" when X = 100 AND Y = 3 else
"010101010101" when X = 101 AND Y = 3 else
"010101010101" when X = 102 AND Y = 3 else
"010101010101" when X = 103 AND Y = 3 else
"010101010101" when X = 104 AND Y = 3 else
"010101010101" when X = 105 AND Y = 3 else
"010101010101" when X = 106 AND Y = 3 else
"010101010101" when X = 107 AND Y = 3 else
"010101010101" when X = 108 AND Y = 3 else
"010101010101" when X = 109 AND Y = 3 else
"010101010101" when X = 110 AND Y = 3 else
"010101010101" when X = 111 AND Y = 3 else
"010101010101" when X = 112 AND Y = 3 else
"010101010101" when X = 113 AND Y = 3 else
"010101010101" when X = 114 AND Y = 3 else
"010101010101" when X = 115 AND Y = 3 else
"010101010101" when X = 116 AND Y = 3 else
"010101010101" when X = 117 AND Y = 3 else
"010101010101" when X = 118 AND Y = 3 else
"010101010101" when X = 119 AND Y = 3 else
"010101010101" when X = 120 AND Y = 3 else
"010101010101" when X = 121 AND Y = 3 else
"010101010101" when X = 122 AND Y = 3 else
"010101010101" when X = 123 AND Y = 3 else
"010101010101" when X = 124 AND Y = 3 else
"010101010101" when X = 125 AND Y = 3 else
"010101010101" when X = 126 AND Y = 3 else
"010101010101" when X = 127 AND Y = 3 else
"010101010101" when X = 128 AND Y = 3 else
"010101010101" when X = 129 AND Y = 3 else
"010101010101" when X = 130 AND Y = 3 else
"010101010101" when X = 131 AND Y = 3 else
"010101010101" when X = 132 AND Y = 3 else
"010101010101" when X = 133 AND Y = 3 else
"010101010101" when X = 134 AND Y = 3 else
"010101010101" when X = 135 AND Y = 3 else
"010101010101" when X = 136 AND Y = 3 else
"010101010101" when X = 137 AND Y = 3 else
"010101010101" when X = 138 AND Y = 3 else
"010101010101" when X = 139 AND Y = 3 else
"010101010101" when X = 140 AND Y = 3 else
"010101010101" when X = 141 AND Y = 3 else
"010101010101" when X = 142 AND Y = 3 else
"010101010101" when X = 143 AND Y = 3 else
"010101010101" when X = 144 AND Y = 3 else
"010101010101" when X = 145 AND Y = 3 else
"010101010101" when X = 146 AND Y = 3 else
"010101010101" when X = 147 AND Y = 3 else
"010101010101" when X = 148 AND Y = 3 else
"010101010101" when X = 149 AND Y = 3 else
"010101010101" when X = 150 AND Y = 3 else
"010101010101" when X = 151 AND Y = 3 else
"010101010101" when X = 152 AND Y = 3 else
"010101010101" when X = 153 AND Y = 3 else
"010101010101" when X = 154 AND Y = 3 else
"010101010101" when X = 155 AND Y = 3 else
"010101010101" when X = 156 AND Y = 3 else
"010101010101" when X = 157 AND Y = 3 else
"010101010101" when X = 158 AND Y = 3 else
"010101010101" when X = 159 AND Y = 3 else
"010101010101" when X = 160 AND Y = 3 else
"010101010101" when X = 161 AND Y = 3 else
"010101010101" when X = 162 AND Y = 3 else
"010101010101" when X = 163 AND Y = 3 else
"010101010101" when X = 164 AND Y = 3 else
"010101010101" when X = 165 AND Y = 3 else
"010101010101" when X = 166 AND Y = 3 else
"010101010101" when X = 167 AND Y = 3 else
"010101010101" when X = 168 AND Y = 3 else
"010101010101" when X = 169 AND Y = 3 else
"010101010101" when X = 170 AND Y = 3 else
"010101010101" when X = 171 AND Y = 3 else
"010101010101" when X = 172 AND Y = 3 else
"010101010101" when X = 173 AND Y = 3 else
"010101010101" when X = 174 AND Y = 3 else
"010101010101" when X = 175 AND Y = 3 else
"010101010101" when X = 176 AND Y = 3 else
"010101010101" when X = 177 AND Y = 3 else
"010101010101" when X = 178 AND Y = 3 else
"010101010101" when X = 179 AND Y = 3 else
"010101010101" when X = 180 AND Y = 3 else
"010101010101" when X = 181 AND Y = 3 else
"010101010101" when X = 182 AND Y = 3 else
"010101010101" when X = 183 AND Y = 3 else
"010101010101" when X = 184 AND Y = 3 else
"010101010101" when X = 185 AND Y = 3 else
"010101010101" when X = 186 AND Y = 3 else
"010101010101" when X = 187 AND Y = 3 else
"010101010101" when X = 188 AND Y = 3 else
"010101010101" when X = 189 AND Y = 3 else
"010101010101" when X = 190 AND Y = 3 else
"010101010101" when X = 191 AND Y = 3 else
"010101010101" when X = 192 AND Y = 3 else
"010101010101" when X = 193 AND Y = 3 else
"010101010101" when X = 194 AND Y = 3 else
"010101010101" when X = 195 AND Y = 3 else
"010101010101" when X = 196 AND Y = 3 else
"010101010101" when X = 197 AND Y = 3 else
"010101010101" when X = 198 AND Y = 3 else
"010101010101" when X = 199 AND Y = 3 else
"010101010101" when X = 200 AND Y = 3 else
"010101010101" when X = 201 AND Y = 3 else
"010101010101" when X = 202 AND Y = 3 else
"010101010101" when X = 203 AND Y = 3 else
"010101010101" when X = 204 AND Y = 3 else
"010101010101" when X = 205 AND Y = 3 else
"010101010101" when X = 206 AND Y = 3 else
"010101010101" when X = 207 AND Y = 3 else
"010101010101" when X = 208 AND Y = 3 else
"010101010101" when X = 209 AND Y = 3 else
"010101010101" when X = 210 AND Y = 3 else
"010101010101" when X = 211 AND Y = 3 else
"010101010101" when X = 212 AND Y = 3 else
"010101010101" when X = 213 AND Y = 3 else
"010101010101" when X = 214 AND Y = 3 else
"010101010101" when X = 215 AND Y = 3 else
"010101010101" when X = 216 AND Y = 3 else
"010101010101" when X = 217 AND Y = 3 else
"010101010101" when X = 218 AND Y = 3 else
"010101010101" when X = 219 AND Y = 3 else
"010101010101" when X = 220 AND Y = 3 else
"010101010101" when X = 221 AND Y = 3 else
"010101010101" when X = 222 AND Y = 3 else
"010101010101" when X = 223 AND Y = 3 else
"010101010101" when X = 224 AND Y = 3 else
"010101010101" when X = 225 AND Y = 3 else
"010101010101" when X = 226 AND Y = 3 else
"111011101110" when X = 227 AND Y = 3 else
"111011101110" when X = 228 AND Y = 3 else
"111011101110" when X = 229 AND Y = 3 else
"111011101110" when X = 230 AND Y = 3 else
"010101010101" when X = 231 AND Y = 3 else
"010101010101" when X = 232 AND Y = 3 else
"010101010101" when X = 233 AND Y = 3 else
"010101010101" when X = 234 AND Y = 3 else
"010101010101" when X = 235 AND Y = 3 else
"010101010101" when X = 236 AND Y = 3 else
"010101010101" when X = 237 AND Y = 3 else
"010101010101" when X = 238 AND Y = 3 else
"010101010101" when X = 239 AND Y = 3 else
"111011101110" when X = 240 AND Y = 3 else
"111011101110" when X = 241 AND Y = 3 else
"111011101110" when X = 242 AND Y = 3 else
"111011101110" when X = 243 AND Y = 3 else
"111011101110" when X = 244 AND Y = 3 else
"111011101110" when X = 245 AND Y = 3 else
"111011101110" when X = 246 AND Y = 3 else
"111011101110" when X = 247 AND Y = 3 else
"111011101110" when X = 248 AND Y = 3 else
"111011101110" when X = 249 AND Y = 3 else
"111011101110" when X = 250 AND Y = 3 else
"111011101110" when X = 251 AND Y = 3 else
"111011101110" when X = 252 AND Y = 3 else
"111011101110" when X = 253 AND Y = 3 else
"111011101110" when X = 254 AND Y = 3 else
"111011101110" when X = 255 AND Y = 3 else
"111000100000" when X = 0 AND Y = 4 else
"111000100000" when X = 1 AND Y = 4 else
"111000100000" when X = 2 AND Y = 4 else
"111000100000" when X = 3 AND Y = 4 else
"111000100000" when X = 4 AND Y = 4 else
"111000100000" when X = 5 AND Y = 4 else
"111000100000" when X = 6 AND Y = 4 else
"111000100000" when X = 7 AND Y = 4 else
"111000100000" when X = 8 AND Y = 4 else
"111000100000" when X = 9 AND Y = 4 else
"111000100000" when X = 10 AND Y = 4 else
"111000100000" when X = 11 AND Y = 4 else
"111000100000" when X = 12 AND Y = 4 else
"111000100000" when X = 13 AND Y = 4 else
"111000100000" when X = 14 AND Y = 4 else
"111000100000" when X = 15 AND Y = 4 else
"010101010101" when X = 16 AND Y = 4 else
"010101010101" when X = 17 AND Y = 4 else
"010101010101" when X = 18 AND Y = 4 else
"010101010101" when X = 19 AND Y = 4 else
"010101010101" when X = 20 AND Y = 4 else
"010101010101" when X = 21 AND Y = 4 else
"010101010101" when X = 22 AND Y = 4 else
"010101010101" when X = 23 AND Y = 4 else
"010101010101" when X = 24 AND Y = 4 else
"111011100000" when X = 25 AND Y = 4 else
"111011100000" when X = 26 AND Y = 4 else
"111011100000" when X = 27 AND Y = 4 else
"111011100000" when X = 28 AND Y = 4 else
"010101010101" when X = 29 AND Y = 4 else
"010101010101" when X = 30 AND Y = 4 else
"010101010101" when X = 31 AND Y = 4 else
"010101010101" when X = 32 AND Y = 4 else
"010101010101" when X = 33 AND Y = 4 else
"010101010101" when X = 34 AND Y = 4 else
"010101010101" when X = 35 AND Y = 4 else
"010101010101" when X = 36 AND Y = 4 else
"010101010101" when X = 37 AND Y = 4 else
"010101010101" when X = 38 AND Y = 4 else
"010101010101" when X = 39 AND Y = 4 else
"010101010101" when X = 40 AND Y = 4 else
"010101010101" when X = 41 AND Y = 4 else
"010101010101" when X = 42 AND Y = 4 else
"010101010101" when X = 43 AND Y = 4 else
"010101010101" when X = 44 AND Y = 4 else
"010101010101" when X = 45 AND Y = 4 else
"010101010101" when X = 46 AND Y = 4 else
"010101010101" when X = 47 AND Y = 4 else
"010101010101" when X = 48 AND Y = 4 else
"010101010101" when X = 49 AND Y = 4 else
"010101010101" when X = 50 AND Y = 4 else
"010101010101" when X = 51 AND Y = 4 else
"010101010101" when X = 52 AND Y = 4 else
"010101010101" when X = 53 AND Y = 4 else
"010101010101" when X = 54 AND Y = 4 else
"010101010101" when X = 55 AND Y = 4 else
"010101010101" when X = 56 AND Y = 4 else
"010101010101" when X = 57 AND Y = 4 else
"010101010101" when X = 58 AND Y = 4 else
"010101010101" when X = 59 AND Y = 4 else
"010101010101" when X = 60 AND Y = 4 else
"010101010101" when X = 61 AND Y = 4 else
"010101010101" when X = 62 AND Y = 4 else
"010101010101" when X = 63 AND Y = 4 else
"010101010101" when X = 64 AND Y = 4 else
"010101010101" when X = 65 AND Y = 4 else
"010101010101" when X = 66 AND Y = 4 else
"010101010101" when X = 67 AND Y = 4 else
"010101010101" when X = 68 AND Y = 4 else
"010101010101" when X = 69 AND Y = 4 else
"010101010101" when X = 70 AND Y = 4 else
"010101010101" when X = 71 AND Y = 4 else
"010101010101" when X = 72 AND Y = 4 else
"010101010101" when X = 73 AND Y = 4 else
"010101010101" when X = 74 AND Y = 4 else
"010101010101" when X = 75 AND Y = 4 else
"010101010101" when X = 76 AND Y = 4 else
"010101010101" when X = 77 AND Y = 4 else
"010101010101" when X = 78 AND Y = 4 else
"010101010101" when X = 79 AND Y = 4 else
"010101010101" when X = 80 AND Y = 4 else
"010101010101" when X = 81 AND Y = 4 else
"010101010101" when X = 82 AND Y = 4 else
"010101010101" when X = 83 AND Y = 4 else
"010101010101" when X = 84 AND Y = 4 else
"010101010101" when X = 85 AND Y = 4 else
"010101010101" when X = 86 AND Y = 4 else
"010101010101" when X = 87 AND Y = 4 else
"010101010101" when X = 88 AND Y = 4 else
"010101010101" when X = 89 AND Y = 4 else
"010101010101" when X = 90 AND Y = 4 else
"010101010101" when X = 91 AND Y = 4 else
"010101010101" when X = 92 AND Y = 4 else
"010101010101" when X = 93 AND Y = 4 else
"010101010101" when X = 94 AND Y = 4 else
"010101010101" when X = 95 AND Y = 4 else
"010101010101" when X = 96 AND Y = 4 else
"010101010101" when X = 97 AND Y = 4 else
"010101010101" when X = 98 AND Y = 4 else
"010101010101" when X = 99 AND Y = 4 else
"010101010101" when X = 100 AND Y = 4 else
"010101010101" when X = 101 AND Y = 4 else
"010101010101" when X = 102 AND Y = 4 else
"010101010101" when X = 103 AND Y = 4 else
"010101010101" when X = 104 AND Y = 4 else
"010101010101" when X = 105 AND Y = 4 else
"010101010101" when X = 106 AND Y = 4 else
"010101010101" when X = 107 AND Y = 4 else
"010101010101" when X = 108 AND Y = 4 else
"010101010101" when X = 109 AND Y = 4 else
"010101010101" when X = 110 AND Y = 4 else
"010101010101" when X = 111 AND Y = 4 else
"010101010101" when X = 112 AND Y = 4 else
"010101010101" when X = 113 AND Y = 4 else
"010101010101" when X = 114 AND Y = 4 else
"010101010101" when X = 115 AND Y = 4 else
"010101010101" when X = 116 AND Y = 4 else
"010101010101" when X = 117 AND Y = 4 else
"010101010101" when X = 118 AND Y = 4 else
"010101010101" when X = 119 AND Y = 4 else
"010101010101" when X = 120 AND Y = 4 else
"010101010101" when X = 121 AND Y = 4 else
"010101010101" when X = 122 AND Y = 4 else
"010101010101" when X = 123 AND Y = 4 else
"010101010101" when X = 124 AND Y = 4 else
"010101010101" when X = 125 AND Y = 4 else
"111011101110" when X = 126 AND Y = 4 else
"111011101110" when X = 127 AND Y = 4 else
"111011101110" when X = 128 AND Y = 4 else
"111011101110" when X = 129 AND Y = 4 else
"010101010101" when X = 130 AND Y = 4 else
"010101010101" when X = 131 AND Y = 4 else
"010101010101" when X = 132 AND Y = 4 else
"010101010101" when X = 133 AND Y = 4 else
"010101010101" when X = 134 AND Y = 4 else
"010101010101" when X = 135 AND Y = 4 else
"010101010101" when X = 136 AND Y = 4 else
"010101010101" when X = 137 AND Y = 4 else
"010101010101" when X = 138 AND Y = 4 else
"010101010101" when X = 139 AND Y = 4 else
"010101010101" when X = 140 AND Y = 4 else
"010101010101" when X = 141 AND Y = 4 else
"010101010101" when X = 142 AND Y = 4 else
"010101010101" when X = 143 AND Y = 4 else
"010101010101" when X = 144 AND Y = 4 else
"010101010101" when X = 145 AND Y = 4 else
"010101010101" when X = 146 AND Y = 4 else
"010101010101" when X = 147 AND Y = 4 else
"010101010101" when X = 148 AND Y = 4 else
"010101010101" when X = 149 AND Y = 4 else
"010101010101" when X = 150 AND Y = 4 else
"010101010101" when X = 151 AND Y = 4 else
"010101010101" when X = 152 AND Y = 4 else
"010101010101" when X = 153 AND Y = 4 else
"010101010101" when X = 154 AND Y = 4 else
"010101010101" when X = 155 AND Y = 4 else
"010101010101" when X = 156 AND Y = 4 else
"010101010101" when X = 157 AND Y = 4 else
"010101010101" when X = 158 AND Y = 4 else
"010101010101" when X = 159 AND Y = 4 else
"010101010101" when X = 160 AND Y = 4 else
"010101010101" when X = 161 AND Y = 4 else
"010101010101" when X = 162 AND Y = 4 else
"010101010101" when X = 163 AND Y = 4 else
"010101010101" when X = 164 AND Y = 4 else
"010101010101" when X = 165 AND Y = 4 else
"010101010101" when X = 166 AND Y = 4 else
"010101010101" when X = 167 AND Y = 4 else
"010101010101" when X = 168 AND Y = 4 else
"010101010101" when X = 169 AND Y = 4 else
"010101010101" when X = 170 AND Y = 4 else
"010101010101" when X = 171 AND Y = 4 else
"010101010101" when X = 172 AND Y = 4 else
"010101010101" when X = 173 AND Y = 4 else
"010101010101" when X = 174 AND Y = 4 else
"010101010101" when X = 175 AND Y = 4 else
"010101010101" when X = 176 AND Y = 4 else
"010101010101" when X = 177 AND Y = 4 else
"010101010101" when X = 178 AND Y = 4 else
"010101010101" when X = 179 AND Y = 4 else
"010101010101" when X = 180 AND Y = 4 else
"010101010101" when X = 181 AND Y = 4 else
"010101010101" when X = 182 AND Y = 4 else
"010101010101" when X = 183 AND Y = 4 else
"010101010101" when X = 184 AND Y = 4 else
"010101010101" when X = 185 AND Y = 4 else
"010101010101" when X = 186 AND Y = 4 else
"010101010101" when X = 187 AND Y = 4 else
"010101010101" when X = 188 AND Y = 4 else
"010101010101" when X = 189 AND Y = 4 else
"010101010101" when X = 190 AND Y = 4 else
"010101010101" when X = 191 AND Y = 4 else
"010101010101" when X = 192 AND Y = 4 else
"010101010101" when X = 193 AND Y = 4 else
"010101010101" when X = 194 AND Y = 4 else
"010101010101" when X = 195 AND Y = 4 else
"010101010101" when X = 196 AND Y = 4 else
"010101010101" when X = 197 AND Y = 4 else
"010101010101" when X = 198 AND Y = 4 else
"010101010101" when X = 199 AND Y = 4 else
"010101010101" when X = 200 AND Y = 4 else
"010101010101" when X = 201 AND Y = 4 else
"010101010101" when X = 202 AND Y = 4 else
"010101010101" when X = 203 AND Y = 4 else
"010101010101" when X = 204 AND Y = 4 else
"010101010101" when X = 205 AND Y = 4 else
"010101010101" when X = 206 AND Y = 4 else
"010101010101" when X = 207 AND Y = 4 else
"010101010101" when X = 208 AND Y = 4 else
"010101010101" when X = 209 AND Y = 4 else
"010101010101" when X = 210 AND Y = 4 else
"010101010101" when X = 211 AND Y = 4 else
"010101010101" when X = 212 AND Y = 4 else
"010101010101" when X = 213 AND Y = 4 else
"010101010101" when X = 214 AND Y = 4 else
"010101010101" when X = 215 AND Y = 4 else
"010101010101" when X = 216 AND Y = 4 else
"010101010101" when X = 217 AND Y = 4 else
"010101010101" when X = 218 AND Y = 4 else
"010101010101" when X = 219 AND Y = 4 else
"010101010101" when X = 220 AND Y = 4 else
"010101010101" when X = 221 AND Y = 4 else
"010101010101" when X = 222 AND Y = 4 else
"010101010101" when X = 223 AND Y = 4 else
"010101010101" when X = 224 AND Y = 4 else
"010101010101" when X = 225 AND Y = 4 else
"010101010101" when X = 226 AND Y = 4 else
"111011100000" when X = 227 AND Y = 4 else
"111011100000" when X = 228 AND Y = 4 else
"111011100000" when X = 229 AND Y = 4 else
"111011100000" when X = 230 AND Y = 4 else
"010101010101" when X = 231 AND Y = 4 else
"010101010101" when X = 232 AND Y = 4 else
"010101010101" when X = 233 AND Y = 4 else
"010101010101" when X = 234 AND Y = 4 else
"010101010101" when X = 235 AND Y = 4 else
"010101010101" when X = 236 AND Y = 4 else
"010101010101" when X = 237 AND Y = 4 else
"010101010101" when X = 238 AND Y = 4 else
"010101010101" when X = 239 AND Y = 4 else
"111000100000" when X = 240 AND Y = 4 else
"111000100000" when X = 241 AND Y = 4 else
"111000100000" when X = 242 AND Y = 4 else
"111000100000" when X = 243 AND Y = 4 else
"111000100000" when X = 244 AND Y = 4 else
"111000100000" when X = 245 AND Y = 4 else
"111000100000" when X = 246 AND Y = 4 else
"111000100000" when X = 247 AND Y = 4 else
"111000100000" when X = 248 AND Y = 4 else
"111000100000" when X = 249 AND Y = 4 else
"111000100000" when X = 250 AND Y = 4 else
"111000100000" when X = 251 AND Y = 4 else
"111000100000" when X = 252 AND Y = 4 else
"111000100000" when X = 253 AND Y = 4 else
"111000100000" when X = 254 AND Y = 4 else
"111000100000" when X = 255 AND Y = 4 else
"111011101110" when X = 0 AND Y = 5 else
"111011101110" when X = 1 AND Y = 5 else
"111011101110" when X = 2 AND Y = 5 else
"111011101110" when X = 3 AND Y = 5 else
"111011101110" when X = 4 AND Y = 5 else
"111011101110" when X = 5 AND Y = 5 else
"111011101110" when X = 6 AND Y = 5 else
"111011101110" when X = 7 AND Y = 5 else
"111011101110" when X = 8 AND Y = 5 else
"111011101110" when X = 9 AND Y = 5 else
"111011101110" when X = 10 AND Y = 5 else
"111011101110" when X = 11 AND Y = 5 else
"111011101110" when X = 12 AND Y = 5 else
"111011101110" when X = 13 AND Y = 5 else
"111011101110" when X = 14 AND Y = 5 else
"111011101110" when X = 15 AND Y = 5 else
"010101010101" when X = 16 AND Y = 5 else
"010101010101" when X = 17 AND Y = 5 else
"010101010101" when X = 18 AND Y = 5 else
"010101010101" when X = 19 AND Y = 5 else
"010101010101" when X = 20 AND Y = 5 else
"010101010101" when X = 21 AND Y = 5 else
"010101010101" when X = 22 AND Y = 5 else
"010101010101" when X = 23 AND Y = 5 else
"010101010101" when X = 24 AND Y = 5 else
"111011100000" when X = 25 AND Y = 5 else
"111011100000" when X = 26 AND Y = 5 else
"111011100000" when X = 27 AND Y = 5 else
"111011100000" when X = 28 AND Y = 5 else
"010101010101" when X = 29 AND Y = 5 else
"010101010101" when X = 30 AND Y = 5 else
"010101010101" when X = 31 AND Y = 5 else
"010101010101" when X = 32 AND Y = 5 else
"010101010101" when X = 33 AND Y = 5 else
"010101010101" when X = 34 AND Y = 5 else
"010101010101" when X = 35 AND Y = 5 else
"010101010101" when X = 36 AND Y = 5 else
"010101010101" when X = 37 AND Y = 5 else
"010101010101" when X = 38 AND Y = 5 else
"010101010101" when X = 39 AND Y = 5 else
"010101010101" when X = 40 AND Y = 5 else
"010101010101" when X = 41 AND Y = 5 else
"010101010101" when X = 42 AND Y = 5 else
"010101010101" when X = 43 AND Y = 5 else
"010101010101" when X = 44 AND Y = 5 else
"010101010101" when X = 45 AND Y = 5 else
"010101010101" when X = 46 AND Y = 5 else
"010101010101" when X = 47 AND Y = 5 else
"010101010101" when X = 48 AND Y = 5 else
"010101010101" when X = 49 AND Y = 5 else
"010101010101" when X = 50 AND Y = 5 else
"010101010101" when X = 51 AND Y = 5 else
"010101010101" when X = 52 AND Y = 5 else
"010101010101" when X = 53 AND Y = 5 else
"010101010101" when X = 54 AND Y = 5 else
"010101010101" when X = 55 AND Y = 5 else
"010101010101" when X = 56 AND Y = 5 else
"010101010101" when X = 57 AND Y = 5 else
"010101010101" when X = 58 AND Y = 5 else
"010101010101" when X = 59 AND Y = 5 else
"010101010101" when X = 60 AND Y = 5 else
"010101010101" when X = 61 AND Y = 5 else
"010101010101" when X = 62 AND Y = 5 else
"010101010101" when X = 63 AND Y = 5 else
"010101010101" when X = 64 AND Y = 5 else
"010101010101" when X = 65 AND Y = 5 else
"010101010101" when X = 66 AND Y = 5 else
"010101010101" when X = 67 AND Y = 5 else
"010101010101" when X = 68 AND Y = 5 else
"010101010101" when X = 69 AND Y = 5 else
"010101010101" when X = 70 AND Y = 5 else
"010101010101" when X = 71 AND Y = 5 else
"010101010101" when X = 72 AND Y = 5 else
"010101010101" when X = 73 AND Y = 5 else
"010101010101" when X = 74 AND Y = 5 else
"010101010101" when X = 75 AND Y = 5 else
"010101010101" when X = 76 AND Y = 5 else
"010101010101" when X = 77 AND Y = 5 else
"010101010101" when X = 78 AND Y = 5 else
"010101010101" when X = 79 AND Y = 5 else
"010101010101" when X = 80 AND Y = 5 else
"010101010101" when X = 81 AND Y = 5 else
"010101010101" when X = 82 AND Y = 5 else
"010101010101" when X = 83 AND Y = 5 else
"010101010101" when X = 84 AND Y = 5 else
"010101010101" when X = 85 AND Y = 5 else
"010101010101" when X = 86 AND Y = 5 else
"010101010101" when X = 87 AND Y = 5 else
"010101010101" when X = 88 AND Y = 5 else
"010101010101" when X = 89 AND Y = 5 else
"010101010101" when X = 90 AND Y = 5 else
"010101010101" when X = 91 AND Y = 5 else
"010101010101" when X = 92 AND Y = 5 else
"010101010101" when X = 93 AND Y = 5 else
"010101010101" when X = 94 AND Y = 5 else
"010101010101" when X = 95 AND Y = 5 else
"010101010101" when X = 96 AND Y = 5 else
"010101010101" when X = 97 AND Y = 5 else
"010101010101" when X = 98 AND Y = 5 else
"010101010101" when X = 99 AND Y = 5 else
"010101010101" when X = 100 AND Y = 5 else
"010101010101" when X = 101 AND Y = 5 else
"010101010101" when X = 102 AND Y = 5 else
"010101010101" when X = 103 AND Y = 5 else
"010101010101" when X = 104 AND Y = 5 else
"010101010101" when X = 105 AND Y = 5 else
"010101010101" when X = 106 AND Y = 5 else
"010101010101" when X = 107 AND Y = 5 else
"010101010101" when X = 108 AND Y = 5 else
"010101010101" when X = 109 AND Y = 5 else
"010101010101" when X = 110 AND Y = 5 else
"010101010101" when X = 111 AND Y = 5 else
"010101010101" when X = 112 AND Y = 5 else
"010101010101" when X = 113 AND Y = 5 else
"010101010101" when X = 114 AND Y = 5 else
"010101010101" when X = 115 AND Y = 5 else
"010101010101" when X = 116 AND Y = 5 else
"010101010101" when X = 117 AND Y = 5 else
"010101010101" when X = 118 AND Y = 5 else
"010101010101" when X = 119 AND Y = 5 else
"010101010101" when X = 120 AND Y = 5 else
"010101010101" when X = 121 AND Y = 5 else
"010101010101" when X = 122 AND Y = 5 else
"010101010101" when X = 123 AND Y = 5 else
"010101010101" when X = 124 AND Y = 5 else
"010101010101" when X = 125 AND Y = 5 else
"111011101110" when X = 126 AND Y = 5 else
"111011101110" when X = 127 AND Y = 5 else
"111011101110" when X = 128 AND Y = 5 else
"111011101110" when X = 129 AND Y = 5 else
"010101010101" when X = 130 AND Y = 5 else
"010101010101" when X = 131 AND Y = 5 else
"010101010101" when X = 132 AND Y = 5 else
"010101010101" when X = 133 AND Y = 5 else
"010101010101" when X = 134 AND Y = 5 else
"010101010101" when X = 135 AND Y = 5 else
"010101010101" when X = 136 AND Y = 5 else
"010101010101" when X = 137 AND Y = 5 else
"010101010101" when X = 138 AND Y = 5 else
"010101010101" when X = 139 AND Y = 5 else
"010101010101" when X = 140 AND Y = 5 else
"010101010101" when X = 141 AND Y = 5 else
"010101010101" when X = 142 AND Y = 5 else
"010101010101" when X = 143 AND Y = 5 else
"010101010101" when X = 144 AND Y = 5 else
"010101010101" when X = 145 AND Y = 5 else
"010101010101" when X = 146 AND Y = 5 else
"010101010101" when X = 147 AND Y = 5 else
"010101010101" when X = 148 AND Y = 5 else
"010101010101" when X = 149 AND Y = 5 else
"010101010101" when X = 150 AND Y = 5 else
"010101010101" when X = 151 AND Y = 5 else
"010101010101" when X = 152 AND Y = 5 else
"010101010101" when X = 153 AND Y = 5 else
"010101010101" when X = 154 AND Y = 5 else
"010101010101" when X = 155 AND Y = 5 else
"010101010101" when X = 156 AND Y = 5 else
"010101010101" when X = 157 AND Y = 5 else
"010101010101" when X = 158 AND Y = 5 else
"010101010101" when X = 159 AND Y = 5 else
"010101010101" when X = 160 AND Y = 5 else
"010101010101" when X = 161 AND Y = 5 else
"010101010101" when X = 162 AND Y = 5 else
"010101010101" when X = 163 AND Y = 5 else
"010101010101" when X = 164 AND Y = 5 else
"010101010101" when X = 165 AND Y = 5 else
"010101010101" when X = 166 AND Y = 5 else
"010101010101" when X = 167 AND Y = 5 else
"010101010101" when X = 168 AND Y = 5 else
"010101010101" when X = 169 AND Y = 5 else
"010101010101" when X = 170 AND Y = 5 else
"010101010101" when X = 171 AND Y = 5 else
"010101010101" when X = 172 AND Y = 5 else
"010101010101" when X = 173 AND Y = 5 else
"010101010101" when X = 174 AND Y = 5 else
"010101010101" when X = 175 AND Y = 5 else
"010101010101" when X = 176 AND Y = 5 else
"010101010101" when X = 177 AND Y = 5 else
"010101010101" when X = 178 AND Y = 5 else
"010101010101" when X = 179 AND Y = 5 else
"010101010101" when X = 180 AND Y = 5 else
"010101010101" when X = 181 AND Y = 5 else
"010101010101" when X = 182 AND Y = 5 else
"010101010101" when X = 183 AND Y = 5 else
"010101010101" when X = 184 AND Y = 5 else
"010101010101" when X = 185 AND Y = 5 else
"010101010101" when X = 186 AND Y = 5 else
"010101010101" when X = 187 AND Y = 5 else
"010101010101" when X = 188 AND Y = 5 else
"010101010101" when X = 189 AND Y = 5 else
"010101010101" when X = 190 AND Y = 5 else
"010101010101" when X = 191 AND Y = 5 else
"010101010101" when X = 192 AND Y = 5 else
"010101010101" when X = 193 AND Y = 5 else
"010101010101" when X = 194 AND Y = 5 else
"010101010101" when X = 195 AND Y = 5 else
"010101010101" when X = 196 AND Y = 5 else
"010101010101" when X = 197 AND Y = 5 else
"010101010101" when X = 198 AND Y = 5 else
"010101010101" when X = 199 AND Y = 5 else
"010101010101" when X = 200 AND Y = 5 else
"010101010101" when X = 201 AND Y = 5 else
"010101010101" when X = 202 AND Y = 5 else
"010101010101" when X = 203 AND Y = 5 else
"010101010101" when X = 204 AND Y = 5 else
"010101010101" when X = 205 AND Y = 5 else
"010101010101" when X = 206 AND Y = 5 else
"010101010101" when X = 207 AND Y = 5 else
"010101010101" when X = 208 AND Y = 5 else
"010101010101" when X = 209 AND Y = 5 else
"010101010101" when X = 210 AND Y = 5 else
"010101010101" when X = 211 AND Y = 5 else
"010101010101" when X = 212 AND Y = 5 else
"010101010101" when X = 213 AND Y = 5 else
"010101010101" when X = 214 AND Y = 5 else
"010101010101" when X = 215 AND Y = 5 else
"010101010101" when X = 216 AND Y = 5 else
"010101010101" when X = 217 AND Y = 5 else
"010101010101" when X = 218 AND Y = 5 else
"010101010101" when X = 219 AND Y = 5 else
"010101010101" when X = 220 AND Y = 5 else
"010101010101" when X = 221 AND Y = 5 else
"010101010101" when X = 222 AND Y = 5 else
"010101010101" when X = 223 AND Y = 5 else
"010101010101" when X = 224 AND Y = 5 else
"010101010101" when X = 225 AND Y = 5 else
"010101010101" when X = 226 AND Y = 5 else
"111011100000" when X = 227 AND Y = 5 else
"111011100000" when X = 228 AND Y = 5 else
"111011100000" when X = 229 AND Y = 5 else
"111011100000" when X = 230 AND Y = 5 else
"010101010101" when X = 231 AND Y = 5 else
"010101010101" when X = 232 AND Y = 5 else
"010101010101" when X = 233 AND Y = 5 else
"010101010101" when X = 234 AND Y = 5 else
"010101010101" when X = 235 AND Y = 5 else
"010101010101" when X = 236 AND Y = 5 else
"010101010101" when X = 237 AND Y = 5 else
"010101010101" when X = 238 AND Y = 5 else
"010101010101" when X = 239 AND Y = 5 else
"111011101110" when X = 240 AND Y = 5 else
"111011101110" when X = 241 AND Y = 5 else
"111011101110" when X = 242 AND Y = 5 else
"111011101110" when X = 243 AND Y = 5 else
"111011101110" when X = 244 AND Y = 5 else
"111011101110" when X = 245 AND Y = 5 else
"111011101110" when X = 246 AND Y = 5 else
"111011101110" when X = 247 AND Y = 5 else
"111011101110" when X = 248 AND Y = 5 else
"111011101110" when X = 249 AND Y = 5 else
"111011101110" when X = 250 AND Y = 5 else
"111011101110" when X = 251 AND Y = 5 else
"111011101110" when X = 252 AND Y = 5 else
"111011101110" when X = 253 AND Y = 5 else
"111011101110" when X = 254 AND Y = 5 else
"111011101110" when X = 255 AND Y = 5 else
"111000100000" when X = 0 AND Y = 6 else
"111000100000" when X = 1 AND Y = 6 else
"111000100000" when X = 2 AND Y = 6 else
"111000100000" when X = 3 AND Y = 6 else
"111000100000" when X = 4 AND Y = 6 else
"111000100000" when X = 5 AND Y = 6 else
"111000100000" when X = 6 AND Y = 6 else
"111000100000" when X = 7 AND Y = 6 else
"111000100000" when X = 8 AND Y = 6 else
"111000100000" when X = 9 AND Y = 6 else
"111000100000" when X = 10 AND Y = 6 else
"111000100000" when X = 11 AND Y = 6 else
"111000100000" when X = 12 AND Y = 6 else
"111000100000" when X = 13 AND Y = 6 else
"111000100000" when X = 14 AND Y = 6 else
"111000100000" when X = 15 AND Y = 6 else
"010101010101" when X = 16 AND Y = 6 else
"010101010101" when X = 17 AND Y = 6 else
"010101010101" when X = 18 AND Y = 6 else
"010101010101" when X = 19 AND Y = 6 else
"010101010101" when X = 20 AND Y = 6 else
"010101010101" when X = 21 AND Y = 6 else
"010101010101" when X = 22 AND Y = 6 else
"010101010101" when X = 23 AND Y = 6 else
"010101010101" when X = 24 AND Y = 6 else
"111011100000" when X = 25 AND Y = 6 else
"111011100000" when X = 26 AND Y = 6 else
"111011100000" when X = 27 AND Y = 6 else
"111011100000" when X = 28 AND Y = 6 else
"010101010101" when X = 29 AND Y = 6 else
"010101010101" when X = 30 AND Y = 6 else
"010101010101" when X = 31 AND Y = 6 else
"010101010101" when X = 32 AND Y = 6 else
"010101010101" when X = 33 AND Y = 6 else
"010101010101" when X = 34 AND Y = 6 else
"010101010101" when X = 35 AND Y = 6 else
"010101010101" when X = 36 AND Y = 6 else
"010101010101" when X = 37 AND Y = 6 else
"010101010101" when X = 38 AND Y = 6 else
"010101010101" when X = 39 AND Y = 6 else
"010101010101" when X = 40 AND Y = 6 else
"010101010101" when X = 41 AND Y = 6 else
"010101010101" when X = 42 AND Y = 6 else
"010101010101" when X = 43 AND Y = 6 else
"010101010101" when X = 44 AND Y = 6 else
"010101010101" when X = 45 AND Y = 6 else
"010101010101" when X = 46 AND Y = 6 else
"010101010101" when X = 47 AND Y = 6 else
"010101010101" when X = 48 AND Y = 6 else
"010101010101" when X = 49 AND Y = 6 else
"010101010101" when X = 50 AND Y = 6 else
"010101010101" when X = 51 AND Y = 6 else
"010101010101" when X = 52 AND Y = 6 else
"010101010101" when X = 53 AND Y = 6 else
"010101010101" when X = 54 AND Y = 6 else
"010101010101" when X = 55 AND Y = 6 else
"010101010101" when X = 56 AND Y = 6 else
"010101010101" when X = 57 AND Y = 6 else
"010101010101" when X = 58 AND Y = 6 else
"010101010101" when X = 59 AND Y = 6 else
"010101010101" when X = 60 AND Y = 6 else
"010101010101" when X = 61 AND Y = 6 else
"010101010101" when X = 62 AND Y = 6 else
"010101010101" when X = 63 AND Y = 6 else
"010101010101" when X = 64 AND Y = 6 else
"010101010101" when X = 65 AND Y = 6 else
"010101010101" when X = 66 AND Y = 6 else
"010101010101" when X = 67 AND Y = 6 else
"010101010101" when X = 68 AND Y = 6 else
"010101010101" when X = 69 AND Y = 6 else
"010101010101" when X = 70 AND Y = 6 else
"010101010101" when X = 71 AND Y = 6 else
"010101010101" when X = 72 AND Y = 6 else
"010101010101" when X = 73 AND Y = 6 else
"010101010101" when X = 74 AND Y = 6 else
"010101010101" when X = 75 AND Y = 6 else
"010101010101" when X = 76 AND Y = 6 else
"010101010101" when X = 77 AND Y = 6 else
"010101010101" when X = 78 AND Y = 6 else
"010101010101" when X = 79 AND Y = 6 else
"010101010101" when X = 80 AND Y = 6 else
"010101010101" when X = 81 AND Y = 6 else
"010101010101" when X = 82 AND Y = 6 else
"010101010101" when X = 83 AND Y = 6 else
"010101010101" when X = 84 AND Y = 6 else
"010101010101" when X = 85 AND Y = 6 else
"010101010101" when X = 86 AND Y = 6 else
"010101010101" when X = 87 AND Y = 6 else
"010101010101" when X = 88 AND Y = 6 else
"010101010101" when X = 89 AND Y = 6 else
"010101010101" when X = 90 AND Y = 6 else
"010101010101" when X = 91 AND Y = 6 else
"010101010101" when X = 92 AND Y = 6 else
"010101010101" when X = 93 AND Y = 6 else
"010101010101" when X = 94 AND Y = 6 else
"010101010101" when X = 95 AND Y = 6 else
"010101010101" when X = 96 AND Y = 6 else
"010101010101" when X = 97 AND Y = 6 else
"010101010101" when X = 98 AND Y = 6 else
"010101010101" when X = 99 AND Y = 6 else
"010101010101" when X = 100 AND Y = 6 else
"010101010101" when X = 101 AND Y = 6 else
"010101010101" when X = 102 AND Y = 6 else
"010101010101" when X = 103 AND Y = 6 else
"010101010101" when X = 104 AND Y = 6 else
"010101010101" when X = 105 AND Y = 6 else
"010101010101" when X = 106 AND Y = 6 else
"010101010101" when X = 107 AND Y = 6 else
"010101010101" when X = 108 AND Y = 6 else
"010101010101" when X = 109 AND Y = 6 else
"010101010101" when X = 110 AND Y = 6 else
"010101010101" when X = 111 AND Y = 6 else
"010101010101" when X = 112 AND Y = 6 else
"010101010101" when X = 113 AND Y = 6 else
"010101010101" when X = 114 AND Y = 6 else
"010101010101" when X = 115 AND Y = 6 else
"010101010101" when X = 116 AND Y = 6 else
"010101010101" when X = 117 AND Y = 6 else
"010101010101" when X = 118 AND Y = 6 else
"010101010101" when X = 119 AND Y = 6 else
"010101010101" when X = 120 AND Y = 6 else
"010101010101" when X = 121 AND Y = 6 else
"010101010101" when X = 122 AND Y = 6 else
"010101010101" when X = 123 AND Y = 6 else
"010101010101" when X = 124 AND Y = 6 else
"010101010101" when X = 125 AND Y = 6 else
"010101010101" when X = 126 AND Y = 6 else
"010101010101" when X = 127 AND Y = 6 else
"010101010101" when X = 128 AND Y = 6 else
"010101010101" when X = 129 AND Y = 6 else
"010101010101" when X = 130 AND Y = 6 else
"010101010101" when X = 131 AND Y = 6 else
"010101010101" when X = 132 AND Y = 6 else
"010101010101" when X = 133 AND Y = 6 else
"010101010101" when X = 134 AND Y = 6 else
"010101010101" when X = 135 AND Y = 6 else
"010101010101" when X = 136 AND Y = 6 else
"010101010101" when X = 137 AND Y = 6 else
"010101010101" when X = 138 AND Y = 6 else
"010101010101" when X = 139 AND Y = 6 else
"010101010101" when X = 140 AND Y = 6 else
"010101010101" when X = 141 AND Y = 6 else
"010101010101" when X = 142 AND Y = 6 else
"010101010101" when X = 143 AND Y = 6 else
"010101010101" when X = 144 AND Y = 6 else
"010101010101" when X = 145 AND Y = 6 else
"010101010101" when X = 146 AND Y = 6 else
"010101010101" when X = 147 AND Y = 6 else
"010101010101" when X = 148 AND Y = 6 else
"010101010101" when X = 149 AND Y = 6 else
"010101010101" when X = 150 AND Y = 6 else
"010101010101" when X = 151 AND Y = 6 else
"010101010101" when X = 152 AND Y = 6 else
"010101010101" when X = 153 AND Y = 6 else
"010101010101" when X = 154 AND Y = 6 else
"010101010101" when X = 155 AND Y = 6 else
"010101010101" when X = 156 AND Y = 6 else
"010101010101" when X = 157 AND Y = 6 else
"010101010101" when X = 158 AND Y = 6 else
"010101010101" when X = 159 AND Y = 6 else
"010101010101" when X = 160 AND Y = 6 else
"010101010101" when X = 161 AND Y = 6 else
"010101010101" when X = 162 AND Y = 6 else
"010101010101" when X = 163 AND Y = 6 else
"010101010101" when X = 164 AND Y = 6 else
"010101010101" when X = 165 AND Y = 6 else
"010101010101" when X = 166 AND Y = 6 else
"010101010101" when X = 167 AND Y = 6 else
"010101010101" when X = 168 AND Y = 6 else
"010101010101" when X = 169 AND Y = 6 else
"010101010101" when X = 170 AND Y = 6 else
"010101010101" when X = 171 AND Y = 6 else
"010101010101" when X = 172 AND Y = 6 else
"010101010101" when X = 173 AND Y = 6 else
"010101010101" when X = 174 AND Y = 6 else
"010101010101" when X = 175 AND Y = 6 else
"010101010101" when X = 176 AND Y = 6 else
"010101010101" when X = 177 AND Y = 6 else
"010101010101" when X = 178 AND Y = 6 else
"010101010101" when X = 179 AND Y = 6 else
"010101010101" when X = 180 AND Y = 6 else
"010101010101" when X = 181 AND Y = 6 else
"010101010101" when X = 182 AND Y = 6 else
"010101010101" when X = 183 AND Y = 6 else
"010101010101" when X = 184 AND Y = 6 else
"010101010101" when X = 185 AND Y = 6 else
"010101010101" when X = 186 AND Y = 6 else
"010101010101" when X = 187 AND Y = 6 else
"010101010101" when X = 188 AND Y = 6 else
"010101010101" when X = 189 AND Y = 6 else
"010101010101" when X = 190 AND Y = 6 else
"010101010101" when X = 191 AND Y = 6 else
"010101010101" when X = 192 AND Y = 6 else
"010101010101" when X = 193 AND Y = 6 else
"010101010101" when X = 194 AND Y = 6 else
"010101010101" when X = 195 AND Y = 6 else
"010101010101" when X = 196 AND Y = 6 else
"010101010101" when X = 197 AND Y = 6 else
"010101010101" when X = 198 AND Y = 6 else
"010101010101" when X = 199 AND Y = 6 else
"010101010101" when X = 200 AND Y = 6 else
"010101010101" when X = 201 AND Y = 6 else
"010101010101" when X = 202 AND Y = 6 else
"010101010101" when X = 203 AND Y = 6 else
"010101010101" when X = 204 AND Y = 6 else
"010101010101" when X = 205 AND Y = 6 else
"010101010101" when X = 206 AND Y = 6 else
"010101010101" when X = 207 AND Y = 6 else
"010101010101" when X = 208 AND Y = 6 else
"010101010101" when X = 209 AND Y = 6 else
"010101010101" when X = 210 AND Y = 6 else
"010101010101" when X = 211 AND Y = 6 else
"010101010101" when X = 212 AND Y = 6 else
"010101010101" when X = 213 AND Y = 6 else
"010101010101" when X = 214 AND Y = 6 else
"010101010101" when X = 215 AND Y = 6 else
"010101010101" when X = 216 AND Y = 6 else
"010101010101" when X = 217 AND Y = 6 else
"010101010101" when X = 218 AND Y = 6 else
"010101010101" when X = 219 AND Y = 6 else
"010101010101" when X = 220 AND Y = 6 else
"010101010101" when X = 221 AND Y = 6 else
"010101010101" when X = 222 AND Y = 6 else
"010101010101" when X = 223 AND Y = 6 else
"010101010101" when X = 224 AND Y = 6 else
"010101010101" when X = 225 AND Y = 6 else
"010101010101" when X = 226 AND Y = 6 else
"111011100000" when X = 227 AND Y = 6 else
"111011100000" when X = 228 AND Y = 6 else
"111011100000" when X = 229 AND Y = 6 else
"111011100000" when X = 230 AND Y = 6 else
"010101010101" when X = 231 AND Y = 6 else
"010101010101" when X = 232 AND Y = 6 else
"010101010101" when X = 233 AND Y = 6 else
"010101010101" when X = 234 AND Y = 6 else
"010101010101" when X = 235 AND Y = 6 else
"010101010101" when X = 236 AND Y = 6 else
"010101010101" when X = 237 AND Y = 6 else
"010101010101" when X = 238 AND Y = 6 else
"010101010101" when X = 239 AND Y = 6 else
"111000100000" when X = 240 AND Y = 6 else
"111000100000" when X = 241 AND Y = 6 else
"111000100000" when X = 242 AND Y = 6 else
"111000100000" when X = 243 AND Y = 6 else
"111000100000" when X = 244 AND Y = 6 else
"111000100000" when X = 245 AND Y = 6 else
"111000100000" when X = 246 AND Y = 6 else
"111000100000" when X = 247 AND Y = 6 else
"111000100000" when X = 248 AND Y = 6 else
"111000100000" when X = 249 AND Y = 6 else
"111000100000" when X = 250 AND Y = 6 else
"111000100000" when X = 251 AND Y = 6 else
"111000100000" when X = 252 AND Y = 6 else
"111000100000" when X = 253 AND Y = 6 else
"111000100000" when X = 254 AND Y = 6 else
"111000100000" when X = 255 AND Y = 6 else
"111011101110" when X = 0 AND Y = 7 else
"111011101110" when X = 1 AND Y = 7 else
"111011101110" when X = 2 AND Y = 7 else
"111011101110" when X = 3 AND Y = 7 else
"111011101110" when X = 4 AND Y = 7 else
"111011101110" when X = 5 AND Y = 7 else
"111011101110" when X = 6 AND Y = 7 else
"111011101110" when X = 7 AND Y = 7 else
"111011101110" when X = 8 AND Y = 7 else
"111011101110" when X = 9 AND Y = 7 else
"111011101110" when X = 10 AND Y = 7 else
"111011101110" when X = 11 AND Y = 7 else
"111011101110" when X = 12 AND Y = 7 else
"111011101110" when X = 13 AND Y = 7 else
"111011101110" when X = 14 AND Y = 7 else
"111011101110" when X = 15 AND Y = 7 else
"010101010101" when X = 16 AND Y = 7 else
"010101010101" when X = 17 AND Y = 7 else
"010101010101" when X = 18 AND Y = 7 else
"010101010101" when X = 19 AND Y = 7 else
"010101010101" when X = 20 AND Y = 7 else
"010101010101" when X = 21 AND Y = 7 else
"010101010101" when X = 22 AND Y = 7 else
"010101010101" when X = 23 AND Y = 7 else
"010101010101" when X = 24 AND Y = 7 else
"111011100000" when X = 25 AND Y = 7 else
"111011100000" when X = 26 AND Y = 7 else
"111011100000" when X = 27 AND Y = 7 else
"111011100000" when X = 28 AND Y = 7 else
"010101010101" when X = 29 AND Y = 7 else
"010101010101" when X = 30 AND Y = 7 else
"010101010101" when X = 31 AND Y = 7 else
"010101010101" when X = 32 AND Y = 7 else
"010101010101" when X = 33 AND Y = 7 else
"010101010101" when X = 34 AND Y = 7 else
"010101010101" when X = 35 AND Y = 7 else
"010101010101" when X = 36 AND Y = 7 else
"010101010101" when X = 37 AND Y = 7 else
"010101010101" when X = 38 AND Y = 7 else
"010101010101" when X = 39 AND Y = 7 else
"010101010101" when X = 40 AND Y = 7 else
"010101010101" when X = 41 AND Y = 7 else
"010101010101" when X = 42 AND Y = 7 else
"010101010101" when X = 43 AND Y = 7 else
"010101010101" when X = 44 AND Y = 7 else
"010101010101" when X = 45 AND Y = 7 else
"010101010101" when X = 46 AND Y = 7 else
"010101010101" when X = 47 AND Y = 7 else
"010101010101" when X = 48 AND Y = 7 else
"010101010101" when X = 49 AND Y = 7 else
"010101010101" when X = 50 AND Y = 7 else
"010101010101" when X = 51 AND Y = 7 else
"010101010101" when X = 52 AND Y = 7 else
"010101010101" when X = 53 AND Y = 7 else
"010101010101" when X = 54 AND Y = 7 else
"010101010101" when X = 55 AND Y = 7 else
"010101010101" when X = 56 AND Y = 7 else
"010101010101" when X = 57 AND Y = 7 else
"010101010101" when X = 58 AND Y = 7 else
"010101010101" when X = 59 AND Y = 7 else
"010101010101" when X = 60 AND Y = 7 else
"010101010101" when X = 61 AND Y = 7 else
"010101010101" when X = 62 AND Y = 7 else
"010101010101" when X = 63 AND Y = 7 else
"010101010101" when X = 64 AND Y = 7 else
"010101010101" when X = 65 AND Y = 7 else
"010101010101" when X = 66 AND Y = 7 else
"010101010101" when X = 67 AND Y = 7 else
"010101010101" when X = 68 AND Y = 7 else
"010101010101" when X = 69 AND Y = 7 else
"010101010101" when X = 70 AND Y = 7 else
"010101010101" when X = 71 AND Y = 7 else
"010101010101" when X = 72 AND Y = 7 else
"010101010101" when X = 73 AND Y = 7 else
"010101010101" when X = 74 AND Y = 7 else
"010101010101" when X = 75 AND Y = 7 else
"010101010101" when X = 76 AND Y = 7 else
"010101010101" when X = 77 AND Y = 7 else
"010101010101" when X = 78 AND Y = 7 else
"010101010101" when X = 79 AND Y = 7 else
"010101010101" when X = 80 AND Y = 7 else
"010101010101" when X = 81 AND Y = 7 else
"010101010101" when X = 82 AND Y = 7 else
"010101010101" when X = 83 AND Y = 7 else
"010101010101" when X = 84 AND Y = 7 else
"010101010101" when X = 85 AND Y = 7 else
"010101010101" when X = 86 AND Y = 7 else
"010101010101" when X = 87 AND Y = 7 else
"010101010101" when X = 88 AND Y = 7 else
"010101010101" when X = 89 AND Y = 7 else
"010101010101" when X = 90 AND Y = 7 else
"010101010101" when X = 91 AND Y = 7 else
"010101010101" when X = 92 AND Y = 7 else
"010101010101" when X = 93 AND Y = 7 else
"010101010101" when X = 94 AND Y = 7 else
"010101010101" when X = 95 AND Y = 7 else
"010101010101" when X = 96 AND Y = 7 else
"010101010101" when X = 97 AND Y = 7 else
"010101010101" when X = 98 AND Y = 7 else
"010101010101" when X = 99 AND Y = 7 else
"010101010101" when X = 100 AND Y = 7 else
"010101010101" when X = 101 AND Y = 7 else
"010101010101" when X = 102 AND Y = 7 else
"010101010101" when X = 103 AND Y = 7 else
"010101010101" when X = 104 AND Y = 7 else
"010101010101" when X = 105 AND Y = 7 else
"010101010101" when X = 106 AND Y = 7 else
"010101010101" when X = 107 AND Y = 7 else
"010101010101" when X = 108 AND Y = 7 else
"010101010101" when X = 109 AND Y = 7 else
"010101010101" when X = 110 AND Y = 7 else
"010101010101" when X = 111 AND Y = 7 else
"010101010101" when X = 112 AND Y = 7 else
"010101010101" when X = 113 AND Y = 7 else
"010101010101" when X = 114 AND Y = 7 else
"010101010101" when X = 115 AND Y = 7 else
"010101010101" when X = 116 AND Y = 7 else
"010101010101" when X = 117 AND Y = 7 else
"010101010101" when X = 118 AND Y = 7 else
"010101010101" when X = 119 AND Y = 7 else
"010101010101" when X = 120 AND Y = 7 else
"010101010101" when X = 121 AND Y = 7 else
"010101010101" when X = 122 AND Y = 7 else
"010101010101" when X = 123 AND Y = 7 else
"010101010101" when X = 124 AND Y = 7 else
"010101010101" when X = 125 AND Y = 7 else
"010101010101" when X = 126 AND Y = 7 else
"010101010101" when X = 127 AND Y = 7 else
"010101010101" when X = 128 AND Y = 7 else
"010101010101" when X = 129 AND Y = 7 else
"010101010101" when X = 130 AND Y = 7 else
"010101010101" when X = 131 AND Y = 7 else
"010101010101" when X = 132 AND Y = 7 else
"010101010101" when X = 133 AND Y = 7 else
"010101010101" when X = 134 AND Y = 7 else
"010101010101" when X = 135 AND Y = 7 else
"010101010101" when X = 136 AND Y = 7 else
"010101010101" when X = 137 AND Y = 7 else
"010101010101" when X = 138 AND Y = 7 else
"010101010101" when X = 139 AND Y = 7 else
"010101010101" when X = 140 AND Y = 7 else
"010101010101" when X = 141 AND Y = 7 else
"010101010101" when X = 142 AND Y = 7 else
"010101010101" when X = 143 AND Y = 7 else
"010101010101" when X = 144 AND Y = 7 else
"010101010101" when X = 145 AND Y = 7 else
"010101010101" when X = 146 AND Y = 7 else
"010101010101" when X = 147 AND Y = 7 else
"010101010101" when X = 148 AND Y = 7 else
"010101010101" when X = 149 AND Y = 7 else
"010101010101" when X = 150 AND Y = 7 else
"010101010101" when X = 151 AND Y = 7 else
"010101010101" when X = 152 AND Y = 7 else
"010101010101" when X = 153 AND Y = 7 else
"010101010101" when X = 154 AND Y = 7 else
"010101010101" when X = 155 AND Y = 7 else
"010101010101" when X = 156 AND Y = 7 else
"010101010101" when X = 157 AND Y = 7 else
"010101010101" when X = 158 AND Y = 7 else
"010101010101" when X = 159 AND Y = 7 else
"010101010101" when X = 160 AND Y = 7 else
"010101010101" when X = 161 AND Y = 7 else
"010101010101" when X = 162 AND Y = 7 else
"010101010101" when X = 163 AND Y = 7 else
"010101010101" when X = 164 AND Y = 7 else
"010101010101" when X = 165 AND Y = 7 else
"010101010101" when X = 166 AND Y = 7 else
"010101010101" when X = 167 AND Y = 7 else
"010101010101" when X = 168 AND Y = 7 else
"010101010101" when X = 169 AND Y = 7 else
"010101010101" when X = 170 AND Y = 7 else
"010101010101" when X = 171 AND Y = 7 else
"010101010101" when X = 172 AND Y = 7 else
"010101010101" when X = 173 AND Y = 7 else
"010101010101" when X = 174 AND Y = 7 else
"010101010101" when X = 175 AND Y = 7 else
"010101010101" when X = 176 AND Y = 7 else
"010101010101" when X = 177 AND Y = 7 else
"010101010101" when X = 178 AND Y = 7 else
"010101010101" when X = 179 AND Y = 7 else
"010101010101" when X = 180 AND Y = 7 else
"010101010101" when X = 181 AND Y = 7 else
"010101010101" when X = 182 AND Y = 7 else
"010101010101" when X = 183 AND Y = 7 else
"010101010101" when X = 184 AND Y = 7 else
"010101010101" when X = 185 AND Y = 7 else
"010101010101" when X = 186 AND Y = 7 else
"010101010101" when X = 187 AND Y = 7 else
"010101010101" when X = 188 AND Y = 7 else
"010101010101" when X = 189 AND Y = 7 else
"010101010101" when X = 190 AND Y = 7 else
"010101010101" when X = 191 AND Y = 7 else
"010101010101" when X = 192 AND Y = 7 else
"010101010101" when X = 193 AND Y = 7 else
"010101010101" when X = 194 AND Y = 7 else
"010101010101" when X = 195 AND Y = 7 else
"010101010101" when X = 196 AND Y = 7 else
"010101010101" when X = 197 AND Y = 7 else
"010101010101" when X = 198 AND Y = 7 else
"010101010101" when X = 199 AND Y = 7 else
"010101010101" when X = 200 AND Y = 7 else
"010101010101" when X = 201 AND Y = 7 else
"010101010101" when X = 202 AND Y = 7 else
"010101010101" when X = 203 AND Y = 7 else
"010101010101" when X = 204 AND Y = 7 else
"010101010101" when X = 205 AND Y = 7 else
"010101010101" when X = 206 AND Y = 7 else
"010101010101" when X = 207 AND Y = 7 else
"010101010101" when X = 208 AND Y = 7 else
"010101010101" when X = 209 AND Y = 7 else
"010101010101" when X = 210 AND Y = 7 else
"010101010101" when X = 211 AND Y = 7 else
"010101010101" when X = 212 AND Y = 7 else
"010101010101" when X = 213 AND Y = 7 else
"010101010101" when X = 214 AND Y = 7 else
"010101010101" when X = 215 AND Y = 7 else
"010101010101" when X = 216 AND Y = 7 else
"010101010101" when X = 217 AND Y = 7 else
"010101010101" when X = 218 AND Y = 7 else
"010101010101" when X = 219 AND Y = 7 else
"010101010101" when X = 220 AND Y = 7 else
"010101010101" when X = 221 AND Y = 7 else
"010101010101" when X = 222 AND Y = 7 else
"010101010101" when X = 223 AND Y = 7 else
"010101010101" when X = 224 AND Y = 7 else
"010101010101" when X = 225 AND Y = 7 else
"010101010101" when X = 226 AND Y = 7 else
"111011100000" when X = 227 AND Y = 7 else
"111011100000" when X = 228 AND Y = 7 else
"111011100000" when X = 229 AND Y = 7 else
"111011100000" when X = 230 AND Y = 7 else
"010101010101" when X = 231 AND Y = 7 else
"010101010101" when X = 232 AND Y = 7 else
"010101010101" when X = 233 AND Y = 7 else
"010101010101" when X = 234 AND Y = 7 else
"010101010101" when X = 235 AND Y = 7 else
"010101010101" when X = 236 AND Y = 7 else
"010101010101" when X = 237 AND Y = 7 else
"010101010101" when X = 238 AND Y = 7 else
"010101010101" when X = 239 AND Y = 7 else
"111011101110" when X = 240 AND Y = 7 else
"111011101110" when X = 241 AND Y = 7 else
"111011101110" when X = 242 AND Y = 7 else
"111011101110" when X = 243 AND Y = 7 else
"111011101110" when X = 244 AND Y = 7 else
"111011101110" when X = 245 AND Y = 7 else
"111011101110" when X = 246 AND Y = 7 else
"111011101110" when X = 247 AND Y = 7 else
"111011101110" when X = 248 AND Y = 7 else
"111011101110" when X = 249 AND Y = 7 else
"111011101110" when X = 250 AND Y = 7 else
"111011101110" when X = 251 AND Y = 7 else
"111011101110" when X = 252 AND Y = 7 else
"111011101110" when X = 253 AND Y = 7 else
"111011101110" when X = 254 AND Y = 7 else
"111011101110" when X = 255 AND Y = 7 else
"000000000000"; -- should never get here
end rtl;
