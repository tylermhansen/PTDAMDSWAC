-- Tyler Hansen
-- CS232 Final Project
-- genSpriteROM.py
-- generates a ROM file in VHDL from a .ppm image

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity cloud is
port(
X	: in INTEGER RANGE 0 TO 1688;
Y	: in INTEGER RANGE 0 TO 1688;
data : out std_logic_vector (12 downto 0)
);

end entity;

architecture rtl of cloud is
begin
data <=
"0000000000000" when X = 0 AND Y = 0 else
"0000000000000" when X = 1 AND Y = 0 else
"0000000000000" when X = 2 AND Y = 0 else
"0000000000000" when X = 3 AND Y = 0 else
"0000000000000" when X = 4 AND Y = 0 else
"0000000000000" when X = 5 AND Y = 0 else
"0000000000000" when X = 6 AND Y = 0 else
"0000000000000" when X = 7 AND Y = 0 else
"0000000000000" when X = 8 AND Y = 0 else
"0000000000000" when X = 9 AND Y = 0 else
"0000000000000" when X = 10 AND Y = 0 else
"0000000000000" when X = 11 AND Y = 0 else
"0000000000000" when X = 12 AND Y = 0 else
"0000000000000" when X = 13 AND Y = 0 else
"0001000100011" when X = 14 AND Y = 0 else
"0011001100111" when X = 15 AND Y = 0 else
"0011001101001" when X = 16 AND Y = 0 else
"0100010001001" when X = 17 AND Y = 0 else
"1100110011001" when X = 18 AND Y = 0 else
"1111111111111" when X = 19 AND Y = 0 else
"1111111111111" when X = 20 AND Y = 0 else
"1111111111111" when X = 21 AND Y = 0 else
"1111111111111" when X = 22 AND Y = 0 else
"1111111111111" when X = 23 AND Y = 0 else
"1111111111111" when X = 24 AND Y = 0 else
"1111111111111" when X = 25 AND Y = 0 else
"1111111111111" when X = 26 AND Y = 0 else
"1111111111111" when X = 27 AND Y = 0 else
"1111111111111" when X = 28 AND Y = 0 else
"1111111111111" when X = 29 AND Y = 0 else
"1111111111111" when X = 30 AND Y = 0 else
"1111111111111" when X = 31 AND Y = 0 else
"1010101010101" when X = 32 AND Y = 0 else
"0010001000101" when X = 33 AND Y = 0 else
"0000000000000" when X = 34 AND Y = 0 else
"0000000000000" when X = 35 AND Y = 0 else
"0000000000000" when X = 36 AND Y = 0 else
"0000000000000" when X = 37 AND Y = 0 else
"0000000000000" when X = 38 AND Y = 0 else
"0000000000000" when X = 39 AND Y = 0 else
"0000000000000" when X = 40 AND Y = 0 else
"0000000000000" when X = 41 AND Y = 0 else
"0000000000000" when X = 42 AND Y = 0 else
"0000000000000" when X = 43 AND Y = 0 else
"0000000000000" when X = 44 AND Y = 0 else
"0000000000000" when X = 45 AND Y = 0 else
"0000000000000" when X = 46 AND Y = 0 else
"0000000000000" when X = 47 AND Y = 0 else
"0000000000000" when X = 48 AND Y = 0 else
"0000000000000" when X = 49 AND Y = 0 else
"0000000000000" when X = 50 AND Y = 0 else
"0000000000000" when X = 51 AND Y = 0 else
"0000000000000" when X = 52 AND Y = 0 else
"0000000000000" when X = 53 AND Y = 0 else
"0000000000000" when X = 54 AND Y = 0 else
"0000000000000" when X = 55 AND Y = 0 else
"0000000000000" when X = 56 AND Y = 0 else
"0000000000000" when X = 57 AND Y = 0 else
"0000000000000" when X = 58 AND Y = 0 else
"0000000000000" when X = 59 AND Y = 0 else
"0000000000000" when X = 60 AND Y = 0 else
"0000000000000" when X = 61 AND Y = 0 else
"0000000000000" when X = 62 AND Y = 0 else
"0000000000000" when X = 63 AND Y = 0 else
"0000000000000" when X = 64 AND Y = 0 else
"0000000000000" when X = 65 AND Y = 0 else
"0000000000000" when X = 66 AND Y = 0 else
"0000000000000" when X = 67 AND Y = 0 else
"0000000000000" when X = 68 AND Y = 0 else
"0000000000000" when X = 69 AND Y = 0 else
"0000000000000" when X = 70 AND Y = 0 else
"0000000000000" when X = 71 AND Y = 0 else
"0000000000000" when X = 72 AND Y = 0 else
"0000000000000" when X = 73 AND Y = 0 else
"0000000000000" when X = 74 AND Y = 0 else
"0000000000000" when X = 0 AND Y = 1 else
"0000000000000" when X = 1 AND Y = 1 else
"0000000000000" when X = 2 AND Y = 1 else
"0000000000000" when X = 3 AND Y = 1 else
"0000000000000" when X = 4 AND Y = 1 else
"0000000000000" when X = 5 AND Y = 1 else
"0000000000000" when X = 6 AND Y = 1 else
"0000000000000" when X = 7 AND Y = 1 else
"0000000000000" when X = 8 AND Y = 1 else
"0000000000000" when X = 9 AND Y = 1 else
"0000000000000" when X = 10 AND Y = 1 else
"0000000000000" when X = 11 AND Y = 1 else
"0000000000000" when X = 12 AND Y = 1 else
"0000000000001" when X = 13 AND Y = 1 else
"0100010001011" when X = 14 AND Y = 1 else
"1011101111001" when X = 15 AND Y = 1 else
"1100110011011" when X = 16 AND Y = 1 else
"1101110111101" when X = 17 AND Y = 1 else
"1111111111111" when X = 18 AND Y = 1 else
"1111111111111" when X = 19 AND Y = 1 else
"1111111111111" when X = 20 AND Y = 1 else
"1111111111111" when X = 21 AND Y = 1 else
"1111111111111" when X = 22 AND Y = 1 else
"1111111111111" when X = 23 AND Y = 1 else
"1111111111111" when X = 24 AND Y = 1 else
"1111111111111" when X = 25 AND Y = 1 else
"1111111111111" when X = 26 AND Y = 1 else
"1111111111111" when X = 27 AND Y = 1 else
"1111111111111" when X = 28 AND Y = 1 else
"1111111111111" when X = 29 AND Y = 1 else
"1111111111111" when X = 30 AND Y = 1 else
"1111111111111" when X = 31 AND Y = 1 else
"1110111011101" when X = 32 AND Y = 1 else
"1010101010101" when X = 33 AND Y = 1 else
"0000000000001" when X = 34 AND Y = 1 else
"0000000000000" when X = 35 AND Y = 1 else
"0000000000000" when X = 36 AND Y = 1 else
"0000000000000" when X = 37 AND Y = 1 else
"0000000000000" when X = 38 AND Y = 1 else
"0000000000000" when X = 39 AND Y = 1 else
"0000000000000" when X = 40 AND Y = 1 else
"0000000000000" when X = 41 AND Y = 1 else
"0000000000000" when X = 42 AND Y = 1 else
"0000000000000" when X = 43 AND Y = 1 else
"0000000000000" when X = 44 AND Y = 1 else
"0000000000000" when X = 45 AND Y = 1 else
"0000000000000" when X = 46 AND Y = 1 else
"0000000000000" when X = 47 AND Y = 1 else
"0000000000000" when X = 48 AND Y = 1 else
"0000000000000" when X = 49 AND Y = 1 else
"0000000000000" when X = 50 AND Y = 1 else
"0000000000000" when X = 51 AND Y = 1 else
"0000000000000" when X = 52 AND Y = 1 else
"0000000000000" when X = 53 AND Y = 1 else
"0000000000000" when X = 54 AND Y = 1 else
"0000000000000" when X = 55 AND Y = 1 else
"0000000000000" when X = 56 AND Y = 1 else
"0000000000000" when X = 57 AND Y = 1 else
"0000000000000" when X = 58 AND Y = 1 else
"0000000000000" when X = 59 AND Y = 1 else
"0000000000000" when X = 60 AND Y = 1 else
"0000000000000" when X = 61 AND Y = 1 else
"0000000000000" when X = 62 AND Y = 1 else
"0000000000000" when X = 63 AND Y = 1 else
"0000000000000" when X = 64 AND Y = 1 else
"0000000000000" when X = 65 AND Y = 1 else
"0000000000000" when X = 66 AND Y = 1 else
"0000000000000" when X = 67 AND Y = 1 else
"0000000000000" when X = 68 AND Y = 1 else
"0000000000000" when X = 69 AND Y = 1 else
"0000000000000" when X = 70 AND Y = 1 else
"0000000000000" when X = 71 AND Y = 1 else
"0000000000000" when X = 72 AND Y = 1 else
"0000000000000" when X = 73 AND Y = 1 else
"0000000000000" when X = 74 AND Y = 1 else
"0000000000000" when X = 0 AND Y = 2 else
"0000000000000" when X = 1 AND Y = 2 else
"0000000000000" when X = 2 AND Y = 2 else
"0000000000000" when X = 3 AND Y = 2 else
"0000000000000" when X = 4 AND Y = 2 else
"0000000000000" when X = 5 AND Y = 2 else
"0000000000000" when X = 6 AND Y = 2 else
"0000000000000" when X = 7 AND Y = 2 else
"0000000000000" when X = 8 AND Y = 2 else
"0000000000000" when X = 9 AND Y = 2 else
"0000000000000" when X = 10 AND Y = 2 else
"0000000000000" when X = 11 AND Y = 2 else
"0000000000000" when X = 12 AND Y = 2 else
"0101010101101" when X = 13 AND Y = 2 else
"1011101111001" when X = 14 AND Y = 2 else
"1101110111101" when X = 15 AND Y = 2 else
"1110111011111" when X = 16 AND Y = 2 else
"1111111111111" when X = 17 AND Y = 2 else
"1111111111111" when X = 18 AND Y = 2 else
"1111111111111" when X = 19 AND Y = 2 else
"1111111111111" when X = 20 AND Y = 2 else
"1111111111111" when X = 21 AND Y = 2 else
"1111111111111" when X = 22 AND Y = 2 else
"1111111111111" when X = 23 AND Y = 2 else
"1111111111111" when X = 24 AND Y = 2 else
"1111111111111" when X = 25 AND Y = 2 else
"1111111111111" when X = 26 AND Y = 2 else
"1111111111111" when X = 27 AND Y = 2 else
"1111111111111" when X = 28 AND Y = 2 else
"1111111111111" when X = 29 AND Y = 2 else
"1111111111111" when X = 30 AND Y = 2 else
"1111111111111" when X = 31 AND Y = 2 else
"1111111111111" when X = 32 AND Y = 2 else
"1110111011101" when X = 33 AND Y = 2 else
"1010101010101" when X = 34 AND Y = 2 else
"0000000000000" when X = 35 AND Y = 2 else
"0000000000000" when X = 36 AND Y = 2 else
"0000000000000" when X = 37 AND Y = 2 else
"0000000000000" when X = 38 AND Y = 2 else
"0000000000000" when X = 39 AND Y = 2 else
"0000000000000" when X = 40 AND Y = 2 else
"0000000000000" when X = 41 AND Y = 2 else
"0000000000000" when X = 42 AND Y = 2 else
"0000000000000" when X = 43 AND Y = 2 else
"0000000000000" when X = 44 AND Y = 2 else
"0000000000000" when X = 45 AND Y = 2 else
"0000000000000" when X = 46 AND Y = 2 else
"0000000000000" when X = 47 AND Y = 2 else
"0000000000000" when X = 48 AND Y = 2 else
"0000000000000" when X = 49 AND Y = 2 else
"0000000000000" when X = 50 AND Y = 2 else
"0000000000000" when X = 51 AND Y = 2 else
"0000000000000" when X = 52 AND Y = 2 else
"0000000000000" when X = 53 AND Y = 2 else
"0000000000000" when X = 54 AND Y = 2 else
"0000000000000" when X = 55 AND Y = 2 else
"0000000000000" when X = 56 AND Y = 2 else
"0000000000000" when X = 57 AND Y = 2 else
"0000000000000" when X = 58 AND Y = 2 else
"0000000000000" when X = 59 AND Y = 2 else
"0000000000000" when X = 60 AND Y = 2 else
"0000000000000" when X = 61 AND Y = 2 else
"0000000000000" when X = 62 AND Y = 2 else
"0000000000000" when X = 63 AND Y = 2 else
"0000000000000" when X = 64 AND Y = 2 else
"0000000000000" when X = 65 AND Y = 2 else
"0000000000000" when X = 66 AND Y = 2 else
"0000000000000" when X = 67 AND Y = 2 else
"0000000000000" when X = 68 AND Y = 2 else
"0000000000000" when X = 69 AND Y = 2 else
"0000000000000" when X = 70 AND Y = 2 else
"0000000000000" when X = 71 AND Y = 2 else
"0000000000000" when X = 72 AND Y = 2 else
"0000000000000" when X = 73 AND Y = 2 else
"0000000000000" when X = 74 AND Y = 2 else
"0000000000000" when X = 0 AND Y = 3 else
"0000000000000" when X = 1 AND Y = 3 else
"0000000000000" when X = 2 AND Y = 3 else
"0000000000000" when X = 3 AND Y = 3 else
"0000000000000" when X = 4 AND Y = 3 else
"0000000000000" when X = 5 AND Y = 3 else
"0000000000000" when X = 6 AND Y = 3 else
"0000000000000" when X = 7 AND Y = 3 else
"0000000000000" when X = 8 AND Y = 3 else
"0000000000000" when X = 9 AND Y = 3 else
"0000000000000" when X = 10 AND Y = 3 else
"0111011110001" when X = 11 AND Y = 3 else
"1010101010111" when X = 12 AND Y = 3 else
"1011101111001" when X = 13 AND Y = 3 else
"1101110111111" when X = 14 AND Y = 3 else
"1110111011111" when X = 15 AND Y = 3 else
"1111111111111" when X = 16 AND Y = 3 else
"1111111111111" when X = 17 AND Y = 3 else
"1111111111111" when X = 18 AND Y = 3 else
"1111111111111" when X = 19 AND Y = 3 else
"1111111111111" when X = 20 AND Y = 3 else
"1111111111111" when X = 21 AND Y = 3 else
"1111111111111" when X = 22 AND Y = 3 else
"1111111111111" when X = 23 AND Y = 3 else
"1111111111111" when X = 24 AND Y = 3 else
"1111111111111" when X = 25 AND Y = 3 else
"1111111111111" when X = 26 AND Y = 3 else
"1111111111111" when X = 27 AND Y = 3 else
"1111111111111" when X = 28 AND Y = 3 else
"1111111111111" when X = 29 AND Y = 3 else
"1111111111111" when X = 30 AND Y = 3 else
"1111111111111" when X = 31 AND Y = 3 else
"1111111111111" when X = 32 AND Y = 3 else
"1111111111111" when X = 33 AND Y = 3 else
"1110111011101" when X = 34 AND Y = 3 else
"1010101010101" when X = 35 AND Y = 3 else
"0010001000101" when X = 36 AND Y = 3 else
"0000000000000" when X = 37 AND Y = 3 else
"0000000000000" when X = 38 AND Y = 3 else
"0000000000000" when X = 39 AND Y = 3 else
"0000000000000" when X = 40 AND Y = 3 else
"0000000000000" when X = 41 AND Y = 3 else
"0000000000000" when X = 42 AND Y = 3 else
"0000000000000" when X = 43 AND Y = 3 else
"0000000000000" when X = 44 AND Y = 3 else
"0000000000000" when X = 45 AND Y = 3 else
"0000000000000" when X = 46 AND Y = 3 else
"0000000000000" when X = 47 AND Y = 3 else
"0000000000000" when X = 48 AND Y = 3 else
"0000000000000" when X = 49 AND Y = 3 else
"0000000000000" when X = 50 AND Y = 3 else
"0000000000000" when X = 51 AND Y = 3 else
"0000000000000" when X = 52 AND Y = 3 else
"0000000000000" when X = 53 AND Y = 3 else
"0000000000000" when X = 54 AND Y = 3 else
"0000000000000" when X = 55 AND Y = 3 else
"0000000000000" when X = 56 AND Y = 3 else
"0000000000000" when X = 57 AND Y = 3 else
"0000000000000" when X = 58 AND Y = 3 else
"0000000000000" when X = 59 AND Y = 3 else
"0000000000000" when X = 60 AND Y = 3 else
"0000000000000" when X = 61 AND Y = 3 else
"0000000000000" when X = 62 AND Y = 3 else
"0000000000000" when X = 63 AND Y = 3 else
"0000000000000" when X = 64 AND Y = 3 else
"0000000000000" when X = 65 AND Y = 3 else
"0000000000000" when X = 66 AND Y = 3 else
"0000000000000" when X = 67 AND Y = 3 else
"0000000000000" when X = 68 AND Y = 3 else
"0000000000000" when X = 69 AND Y = 3 else
"0000000000000" when X = 70 AND Y = 3 else
"0000000000000" when X = 71 AND Y = 3 else
"0000000000000" when X = 72 AND Y = 3 else
"0000000000000" when X = 73 AND Y = 3 else
"0000000000000" when X = 74 AND Y = 3 else
"0000000000000" when X = 0 AND Y = 4 else
"0000000000000" when X = 1 AND Y = 4 else
"0000000000000" when X = 2 AND Y = 4 else
"0000000000000" when X = 3 AND Y = 4 else
"0000000000000" when X = 4 AND Y = 4 else
"0000000000000" when X = 5 AND Y = 4 else
"0000000000000" when X = 6 AND Y = 4 else
"0000000000000" when X = 7 AND Y = 4 else
"0000000000000" when X = 8 AND Y = 4 else
"0000000000000" when X = 9 AND Y = 4 else
"0100010001111" when X = 10 AND Y = 4 else
"1001101011001" when X = 11 AND Y = 4 else
"1101110111111" when X = 12 AND Y = 4 else
"1101110111111" when X = 13 AND Y = 4 else
"1110111011111" when X = 14 AND Y = 4 else
"1111111111111" when X = 15 AND Y = 4 else
"1111111111111" when X = 16 AND Y = 4 else
"1111111111111" when X = 17 AND Y = 4 else
"1111111111111" when X = 18 AND Y = 4 else
"1111111111111" when X = 19 AND Y = 4 else
"1111111111111" when X = 20 AND Y = 4 else
"1111111111111" when X = 21 AND Y = 4 else
"1111111111111" when X = 22 AND Y = 4 else
"1111111111111" when X = 23 AND Y = 4 else
"1111111111111" when X = 24 AND Y = 4 else
"1111111111111" when X = 25 AND Y = 4 else
"1111111111111" when X = 26 AND Y = 4 else
"1111111111111" when X = 27 AND Y = 4 else
"1111111111111" when X = 28 AND Y = 4 else
"1111111111111" when X = 29 AND Y = 4 else
"1111111111111" when X = 30 AND Y = 4 else
"1111111111111" when X = 31 AND Y = 4 else
"1111111111111" when X = 32 AND Y = 4 else
"1111111111111" when X = 33 AND Y = 4 else
"1111111111111" when X = 34 AND Y = 4 else
"1101110111011" when X = 35 AND Y = 4 else
"0001000100011" when X = 36 AND Y = 4 else
"0000000000000" when X = 37 AND Y = 4 else
"0000000000000" when X = 38 AND Y = 4 else
"0000000000000" when X = 39 AND Y = 4 else
"0000000000000" when X = 40 AND Y = 4 else
"0000000000000" when X = 41 AND Y = 4 else
"0000000000000" when X = 42 AND Y = 4 else
"0000000000000" when X = 43 AND Y = 4 else
"0000000000000" when X = 44 AND Y = 4 else
"0000000000000" when X = 45 AND Y = 4 else
"0000000000000" when X = 46 AND Y = 4 else
"0000000000000" when X = 47 AND Y = 4 else
"0000000000000" when X = 48 AND Y = 4 else
"0000000000000" when X = 49 AND Y = 4 else
"0000000000000" when X = 50 AND Y = 4 else
"0000000000000" when X = 51 AND Y = 4 else
"0000000000000" when X = 52 AND Y = 4 else
"0000000000000" when X = 53 AND Y = 4 else
"0000000000000" when X = 54 AND Y = 4 else
"0000000000000" when X = 55 AND Y = 4 else
"0000000000000" when X = 56 AND Y = 4 else
"0000000000000" when X = 57 AND Y = 4 else
"0000000000000" when X = 58 AND Y = 4 else
"0000000000000" when X = 59 AND Y = 4 else
"0000000000000" when X = 60 AND Y = 4 else
"0000000000000" when X = 61 AND Y = 4 else
"0000000000000" when X = 62 AND Y = 4 else
"0000000000000" when X = 63 AND Y = 4 else
"0000000000000" when X = 64 AND Y = 4 else
"0000000000000" when X = 65 AND Y = 4 else
"0000000000000" when X = 66 AND Y = 4 else
"0000000000000" when X = 67 AND Y = 4 else
"0000000000000" when X = 68 AND Y = 4 else
"0000000000000" when X = 69 AND Y = 4 else
"0000000000000" when X = 70 AND Y = 4 else
"0000000000000" when X = 71 AND Y = 4 else
"0000000000000" when X = 72 AND Y = 4 else
"0000000000000" when X = 73 AND Y = 4 else
"0000000000000" when X = 74 AND Y = 4 else
"0000000000000" when X = 0 AND Y = 5 else
"0000000000000" when X = 1 AND Y = 5 else
"0000000000000" when X = 2 AND Y = 5 else
"0000000000000" when X = 3 AND Y = 5 else
"0000000000000" when X = 4 AND Y = 5 else
"0000000000000" when X = 5 AND Y = 5 else
"0000000000000" when X = 6 AND Y = 5 else
"0000000000000" when X = 7 AND Y = 5 else
"0000000000000" when X = 8 AND Y = 5 else
"0000000000000" when X = 9 AND Y = 5 else
"0110011110101" when X = 10 AND Y = 5 else
"1010101111101" when X = 11 AND Y = 5 else
"1101110111111" when X = 12 AND Y = 5 else
"1101111011111" when X = 13 AND Y = 5 else
"1111111111111" when X = 14 AND Y = 5 else
"1111111111111" when X = 15 AND Y = 5 else
"1111111111111" when X = 16 AND Y = 5 else
"1111111111111" when X = 17 AND Y = 5 else
"1111111111111" when X = 18 AND Y = 5 else
"1111111111111" when X = 19 AND Y = 5 else
"1111111111111" when X = 20 AND Y = 5 else
"1111111111111" when X = 21 AND Y = 5 else
"1111111111111" when X = 22 AND Y = 5 else
"1111111111111" when X = 23 AND Y = 5 else
"1111111111111" when X = 24 AND Y = 5 else
"1111111111111" when X = 25 AND Y = 5 else
"1111111111111" when X = 26 AND Y = 5 else
"1111111111111" when X = 27 AND Y = 5 else
"1111111111111" when X = 28 AND Y = 5 else
"1111111111111" when X = 29 AND Y = 5 else
"1111111111111" when X = 30 AND Y = 5 else
"1111111111111" when X = 31 AND Y = 5 else
"1111111111111" when X = 32 AND Y = 5 else
"1111111111111" when X = 33 AND Y = 5 else
"1111111111111" when X = 34 AND Y = 5 else
"1110111011101" when X = 35 AND Y = 5 else
"1000100010001" when X = 36 AND Y = 5 else
"0001000100011" when X = 37 AND Y = 5 else
"0000000000000" when X = 38 AND Y = 5 else
"0000000000000" when X = 39 AND Y = 5 else
"0000000000000" when X = 40 AND Y = 5 else
"0000000000000" when X = 41 AND Y = 5 else
"0000000000000" when X = 42 AND Y = 5 else
"0000000000000" when X = 43 AND Y = 5 else
"0000000000000" when X = 44 AND Y = 5 else
"0000000000000" when X = 45 AND Y = 5 else
"0000000000000" when X = 46 AND Y = 5 else
"0000000000000" when X = 47 AND Y = 5 else
"0000000000000" when X = 48 AND Y = 5 else
"0000000000000" when X = 49 AND Y = 5 else
"0000000000000" when X = 50 AND Y = 5 else
"0000000000000" when X = 51 AND Y = 5 else
"0000000000000" when X = 52 AND Y = 5 else
"0000000000000" when X = 53 AND Y = 5 else
"0111011101111" when X = 54 AND Y = 5 else
"1001100110011" when X = 55 AND Y = 5 else
"1001100110011" when X = 56 AND Y = 5 else
"1000100010011" when X = 57 AND Y = 5 else
"0111011110001" when X = 58 AND Y = 5 else
"0111011110001" when X = 59 AND Y = 5 else
"0111011110001" when X = 60 AND Y = 5 else
"0111011110001" when X = 61 AND Y = 5 else
"0100010001011" when X = 62 AND Y = 5 else
"0000000000000" when X = 63 AND Y = 5 else
"0000000000000" when X = 64 AND Y = 5 else
"0000000000000" when X = 65 AND Y = 5 else
"0000000000000" when X = 66 AND Y = 5 else
"0000000000000" when X = 67 AND Y = 5 else
"0000000000000" when X = 68 AND Y = 5 else
"0000000000000" when X = 69 AND Y = 5 else
"0000000000000" when X = 70 AND Y = 5 else
"0000000000000" when X = 71 AND Y = 5 else
"0000000000000" when X = 72 AND Y = 5 else
"0000000000000" when X = 73 AND Y = 5 else
"0000000000000" when X = 74 AND Y = 5 else
"0000000000000" when X = 0 AND Y = 6 else
"0000000000000" when X = 1 AND Y = 6 else
"0000000000000" when X = 2 AND Y = 6 else
"0000000000000" when X = 3 AND Y = 6 else
"0000000000000" when X = 4 AND Y = 6 else
"0000000000000" when X = 5 AND Y = 6 else
"0000000000000" when X = 6 AND Y = 6 else
"0000000000000" when X = 7 AND Y = 6 else
"0000000000000" when X = 8 AND Y = 6 else
"0000000000000" when X = 9 AND Y = 6 else
"0110011110101" when X = 10 AND Y = 6 else
"1010101111101" when X = 11 AND Y = 6 else
"1101110111111" when X = 12 AND Y = 6 else
"1101111011111" when X = 13 AND Y = 6 else
"1111111111111" when X = 14 AND Y = 6 else
"1111111111111" when X = 15 AND Y = 6 else
"1111111111111" when X = 16 AND Y = 6 else
"1111111111111" when X = 17 AND Y = 6 else
"1111111111111" when X = 18 AND Y = 6 else
"1111111111111" when X = 19 AND Y = 6 else
"1111111111111" when X = 20 AND Y = 6 else
"1111111111111" when X = 21 AND Y = 6 else
"1111111111111" when X = 22 AND Y = 6 else
"1111111111111" when X = 23 AND Y = 6 else
"1111111111111" when X = 24 AND Y = 6 else
"1111111111111" when X = 25 AND Y = 6 else
"1111111111111" when X = 26 AND Y = 6 else
"1111111111111" when X = 27 AND Y = 6 else
"1111111111111" when X = 28 AND Y = 6 else
"1111111111111" when X = 29 AND Y = 6 else
"1111111111111" when X = 30 AND Y = 6 else
"1111111111111" when X = 31 AND Y = 6 else
"1111111111111" when X = 32 AND Y = 6 else
"1111111111111" when X = 33 AND Y = 6 else
"1111111111111" when X = 34 AND Y = 6 else
"1111111111111" when X = 35 AND Y = 6 else
"1110111011101" when X = 36 AND Y = 6 else
"1000100010001" when X = 37 AND Y = 6 else
"0111011101111" when X = 38 AND Y = 6 else
"0111011101111" when X = 39 AND Y = 6 else
"0111011101111" when X = 40 AND Y = 6 else
"0111011101111" when X = 41 AND Y = 6 else
"0111011101111" when X = 42 AND Y = 6 else
"0110011001101" when X = 43 AND Y = 6 else
"0000000000001" when X = 44 AND Y = 6 else
"0000000000000" when X = 45 AND Y = 6 else
"0000000000000" when X = 46 AND Y = 6 else
"0000000000000" when X = 47 AND Y = 6 else
"0000000000000" when X = 48 AND Y = 6 else
"0000000000000" when X = 49 AND Y = 6 else
"0000000000000" when X = 50 AND Y = 6 else
"0010001000101" when X = 51 AND Y = 6 else
"0111011101111" when X = 52 AND Y = 6 else
"0111011101111" when X = 53 AND Y = 6 else
"1110111011101" when X = 54 AND Y = 6 else
"1111111111111" when X = 55 AND Y = 6 else
"1111111111111" when X = 56 AND Y = 6 else
"1111111111111" when X = 57 AND Y = 6 else
"1101110111111" when X = 58 AND Y = 6 else
"1101110111101" when X = 59 AND Y = 6 else
"1101110111101" when X = 60 AND Y = 6 else
"1101110111101" when X = 61 AND Y = 6 else
"1001100110101" when X = 62 AND Y = 6 else
"0100010001001" when X = 63 AND Y = 6 else
"0000000000000" when X = 64 AND Y = 6 else
"0000000000000" when X = 65 AND Y = 6 else
"0000000000000" when X = 66 AND Y = 6 else
"0000000000000" when X = 67 AND Y = 6 else
"0000000000000" when X = 68 AND Y = 6 else
"0000000000000" when X = 69 AND Y = 6 else
"0000000000000" when X = 70 AND Y = 6 else
"0000000000000" when X = 71 AND Y = 6 else
"0000000000000" when X = 72 AND Y = 6 else
"0000000000000" when X = 73 AND Y = 6 else
"0000000000000" when X = 74 AND Y = 6 else
"0000000000000" when X = 0 AND Y = 7 else
"0000000000000" when X = 1 AND Y = 7 else
"0000000000000" when X = 2 AND Y = 7 else
"0000000000000" when X = 3 AND Y = 7 else
"0000000000000" when X = 4 AND Y = 7 else
"0000000000000" when X = 5 AND Y = 7 else
"0000000000000" when X = 6 AND Y = 7 else
"0000000000000" when X = 7 AND Y = 7 else
"0000000000000" when X = 8 AND Y = 7 else
"0000000000000" when X = 9 AND Y = 7 else
"0110011110101" when X = 10 AND Y = 7 else
"1010101111101" when X = 11 AND Y = 7 else
"1101110111111" when X = 12 AND Y = 7 else
"1101111011111" when X = 13 AND Y = 7 else
"1111111111111" when X = 14 AND Y = 7 else
"1111111111111" when X = 15 AND Y = 7 else
"1111111111111" when X = 16 AND Y = 7 else
"1111111111111" when X = 17 AND Y = 7 else
"1111111111111" when X = 18 AND Y = 7 else
"1111111111111" when X = 19 AND Y = 7 else
"1111111111111" when X = 20 AND Y = 7 else
"1111111111111" when X = 21 AND Y = 7 else
"1111111111111" when X = 22 AND Y = 7 else
"1111111111111" when X = 23 AND Y = 7 else
"1111111111111" when X = 24 AND Y = 7 else
"1111111111111" when X = 25 AND Y = 7 else
"1111111111111" when X = 26 AND Y = 7 else
"1111111111111" when X = 27 AND Y = 7 else
"1111111111111" when X = 28 AND Y = 7 else
"1111111111111" when X = 29 AND Y = 7 else
"1111111111111" when X = 30 AND Y = 7 else
"1111111111111" when X = 31 AND Y = 7 else
"1111111111111" when X = 32 AND Y = 7 else
"1111111111111" when X = 33 AND Y = 7 else
"1111111111111" when X = 34 AND Y = 7 else
"1111111111111" when X = 35 AND Y = 7 else
"1111111111111" when X = 36 AND Y = 7 else
"1111111111111" when X = 37 AND Y = 7 else
"1111111111111" when X = 38 AND Y = 7 else
"1111111111111" when X = 39 AND Y = 7 else
"1111111111111" when X = 40 AND Y = 7 else
"1111111111111" when X = 41 AND Y = 7 else
"1111111111111" when X = 42 AND Y = 7 else
"1110111011101" when X = 43 AND Y = 7 else
"0110011001101" when X = 44 AND Y = 7 else
"0101010101011" when X = 45 AND Y = 7 else
"0010001000101" when X = 46 AND Y = 7 else
"0000000000000" when X = 47 AND Y = 7 else
"0000000000000" when X = 48 AND Y = 7 else
"0011001100111" when X = 49 AND Y = 7 else
"0101010101011" when X = 50 AND Y = 7 else
"1000100010001" when X = 51 AND Y = 7 else
"1110111011101" when X = 52 AND Y = 7 else
"1111111111111" when X = 53 AND Y = 7 else
"1111111111111" when X = 54 AND Y = 7 else
"1111111111111" when X = 55 AND Y = 7 else
"1111111111111" when X = 56 AND Y = 7 else
"1111111111111" when X = 57 AND Y = 7 else
"1111111111111" when X = 58 AND Y = 7 else
"1101111011111" when X = 59 AND Y = 7 else
"1101110111111" when X = 60 AND Y = 7 else
"1101110111111" when X = 61 AND Y = 7 else
"1101110111101" when X = 62 AND Y = 7 else
"1001100110101" when X = 63 AND Y = 7 else
"0011001101001" when X = 64 AND Y = 7 else
"0000000000000" when X = 65 AND Y = 7 else
"0000000000000" when X = 66 AND Y = 7 else
"0000000000000" when X = 67 AND Y = 7 else
"0000000000000" when X = 68 AND Y = 7 else
"0000000000000" when X = 69 AND Y = 7 else
"0000000000000" when X = 70 AND Y = 7 else
"0000000000000" when X = 71 AND Y = 7 else
"0000000000000" when X = 72 AND Y = 7 else
"0000000000000" when X = 73 AND Y = 7 else
"0000000000000" when X = 74 AND Y = 7 else
"0000000000000" when X = 0 AND Y = 8 else
"0000000000000" when X = 1 AND Y = 8 else
"0000000000000" when X = 2 AND Y = 8 else
"0000000000000" when X = 3 AND Y = 8 else
"0000000000000" when X = 4 AND Y = 8 else
"0000000000000" when X = 5 AND Y = 8 else
"0000000000000" when X = 6 AND Y = 8 else
"0000000000000" when X = 7 AND Y = 8 else
"0000000000000" when X = 8 AND Y = 8 else
"0000000000000" when X = 9 AND Y = 8 else
"0110011110101" when X = 10 AND Y = 8 else
"1010101111101" when X = 11 AND Y = 8 else
"1101110111111" when X = 12 AND Y = 8 else
"1101111011111" when X = 13 AND Y = 8 else
"1111111111111" when X = 14 AND Y = 8 else
"1111111111111" when X = 15 AND Y = 8 else
"1111111111111" when X = 16 AND Y = 8 else
"1111111111111" when X = 17 AND Y = 8 else
"1111111111111" when X = 18 AND Y = 8 else
"1111111111111" when X = 19 AND Y = 8 else
"1111111111111" when X = 20 AND Y = 8 else
"1111111111111" when X = 21 AND Y = 8 else
"1111111111111" when X = 22 AND Y = 8 else
"1111111111111" when X = 23 AND Y = 8 else
"1111111111111" when X = 24 AND Y = 8 else
"1111111111111" when X = 25 AND Y = 8 else
"1111111111111" when X = 26 AND Y = 8 else
"1111111111111" when X = 27 AND Y = 8 else
"1111111111111" when X = 28 AND Y = 8 else
"1111111111111" when X = 29 AND Y = 8 else
"1111111111111" when X = 30 AND Y = 8 else
"1111111111111" when X = 31 AND Y = 8 else
"1111111111111" when X = 32 AND Y = 8 else
"1111111111111" when X = 33 AND Y = 8 else
"1111111111111" when X = 34 AND Y = 8 else
"1111111111111" when X = 35 AND Y = 8 else
"1111111111111" when X = 36 AND Y = 8 else
"1111111111111" when X = 37 AND Y = 8 else
"1111111111111" when X = 38 AND Y = 8 else
"1111111111111" when X = 39 AND Y = 8 else
"1111111111111" when X = 40 AND Y = 8 else
"1111111111111" when X = 41 AND Y = 8 else
"1111111111111" when X = 42 AND Y = 8 else
"1111111111111" when X = 43 AND Y = 8 else
"1110111011101" when X = 44 AND Y = 8 else
"1110111011101" when X = 45 AND Y = 8 else
"1000100010001" when X = 46 AND Y = 8 else
"0011001100111" when X = 47 AND Y = 8 else
"0011001100111" when X = 48 AND Y = 8 else
"1010101010101" when X = 49 AND Y = 8 else
"1110111011101" when X = 50 AND Y = 8 else
"1111111111111" when X = 51 AND Y = 8 else
"1111111111111" when X = 52 AND Y = 8 else
"1111111111111" when X = 53 AND Y = 8 else
"1111111111111" when X = 54 AND Y = 8 else
"1111111111111" when X = 55 AND Y = 8 else
"1111111111111" when X = 56 AND Y = 8 else
"1111111111111" when X = 57 AND Y = 8 else
"1111111111111" when X = 58 AND Y = 8 else
"1111111111111" when X = 59 AND Y = 8 else
"1101111011111" when X = 60 AND Y = 8 else
"1101110111111" when X = 61 AND Y = 8 else
"1101110111111" when X = 62 AND Y = 8 else
"1100110111101" when X = 63 AND Y = 8 else
"1001101010111" when X = 64 AND Y = 8 else
"0000000000000" when X = 65 AND Y = 8 else
"0000000000000" when X = 66 AND Y = 8 else
"0000000000000" when X = 67 AND Y = 8 else
"0000000000000" when X = 68 AND Y = 8 else
"0000000000000" when X = 69 AND Y = 8 else
"0000000000000" when X = 70 AND Y = 8 else
"0000000000000" when X = 71 AND Y = 8 else
"0000000000000" when X = 72 AND Y = 8 else
"0000000000000" when X = 73 AND Y = 8 else
"0000000000000" when X = 74 AND Y = 8 else
"0000000000000" when X = 0 AND Y = 9 else
"0000000000000" when X = 1 AND Y = 9 else
"0000000000000" when X = 2 AND Y = 9 else
"0000000000000" when X = 3 AND Y = 9 else
"0000000000000" when X = 4 AND Y = 9 else
"0000000000000" when X = 5 AND Y = 9 else
"0000000000000" when X = 6 AND Y = 9 else
"0000000000000" when X = 7 AND Y = 9 else
"0000000000000" when X = 8 AND Y = 9 else
"0000000000000" when X = 9 AND Y = 9 else
"0110011110101" when X = 10 AND Y = 9 else
"1010101111101" when X = 11 AND Y = 9 else
"1101110111111" when X = 12 AND Y = 9 else
"1101111011111" when X = 13 AND Y = 9 else
"1111111111111" when X = 14 AND Y = 9 else
"1111111111111" when X = 15 AND Y = 9 else
"1111111111111" when X = 16 AND Y = 9 else
"1111111111111" when X = 17 AND Y = 9 else
"1111111111111" when X = 18 AND Y = 9 else
"1111111111111" when X = 19 AND Y = 9 else
"1111111111111" when X = 20 AND Y = 9 else
"1111111111111" when X = 21 AND Y = 9 else
"1111111111111" when X = 22 AND Y = 9 else
"1111111111111" when X = 23 AND Y = 9 else
"1111111111111" when X = 24 AND Y = 9 else
"1111111111111" when X = 25 AND Y = 9 else
"1111111111111" when X = 26 AND Y = 9 else
"1111111111111" when X = 27 AND Y = 9 else
"1111111111111" when X = 28 AND Y = 9 else
"1111111111111" when X = 29 AND Y = 9 else
"1111111111111" when X = 30 AND Y = 9 else
"1111111111111" when X = 31 AND Y = 9 else
"1111111111111" when X = 32 AND Y = 9 else
"1111111111111" when X = 33 AND Y = 9 else
"1111111111111" when X = 34 AND Y = 9 else
"1111111111111" when X = 35 AND Y = 9 else
"1111111111111" when X = 36 AND Y = 9 else
"1111111111111" when X = 37 AND Y = 9 else
"1111111111111" when X = 38 AND Y = 9 else
"1111111111111" when X = 39 AND Y = 9 else
"1111111111111" when X = 40 AND Y = 9 else
"1111111111111" when X = 41 AND Y = 9 else
"1111111111111" when X = 42 AND Y = 9 else
"1111111111111" when X = 43 AND Y = 9 else
"1111111111111" when X = 44 AND Y = 9 else
"1111111111111" when X = 45 AND Y = 9 else
"1110111011101" when X = 46 AND Y = 9 else
"1110111011101" when X = 47 AND Y = 9 else
"1110111011101" when X = 48 AND Y = 9 else
"1110111011101" when X = 49 AND Y = 9 else
"1111111111111" when X = 50 AND Y = 9 else
"1111111111111" when X = 51 AND Y = 9 else
"1111111111111" when X = 52 AND Y = 9 else
"1111111111111" when X = 53 AND Y = 9 else
"1111111111111" when X = 54 AND Y = 9 else
"1111111111111" when X = 55 AND Y = 9 else
"1111111111111" when X = 56 AND Y = 9 else
"1111111111111" when X = 57 AND Y = 9 else
"1111111111111" when X = 58 AND Y = 9 else
"1111111111111" when X = 59 AND Y = 9 else
"1111111111111" when X = 60 AND Y = 9 else
"1101111011111" when X = 61 AND Y = 9 else
"1101110111111" when X = 62 AND Y = 9 else
"1101110111111" when X = 63 AND Y = 9 else
"1010101011001" when X = 64 AND Y = 9 else
"0000000000000" when X = 65 AND Y = 9 else
"0000000000000" when X = 66 AND Y = 9 else
"0000000000000" when X = 67 AND Y = 9 else
"0000000000000" when X = 68 AND Y = 9 else
"0000000000000" when X = 69 AND Y = 9 else
"0000000000000" when X = 70 AND Y = 9 else
"0000000000000" when X = 71 AND Y = 9 else
"0000000000000" when X = 72 AND Y = 9 else
"0000000000000" when X = 73 AND Y = 9 else
"0000000000000" when X = 74 AND Y = 9 else
"0000000000000" when X = 0 AND Y = 10 else
"0000000000000" when X = 1 AND Y = 10 else
"0000000000000" when X = 2 AND Y = 10 else
"0000000000000" when X = 3 AND Y = 10 else
"0000000000000" when X = 4 AND Y = 10 else
"0000000000000" when X = 5 AND Y = 10 else
"0000000000000" when X = 6 AND Y = 10 else
"0000000000000" when X = 7 AND Y = 10 else
"0000000000000" when X = 8 AND Y = 10 else
"0000000000000" when X = 9 AND Y = 10 else
"0110011110101" when X = 10 AND Y = 10 else
"1010101111101" when X = 11 AND Y = 10 else
"1101110111111" when X = 12 AND Y = 10 else
"1101111011111" when X = 13 AND Y = 10 else
"1111111111111" when X = 14 AND Y = 10 else
"1111111111111" when X = 15 AND Y = 10 else
"1111111111111" when X = 16 AND Y = 10 else
"1111111111111" when X = 17 AND Y = 10 else
"1111111111111" when X = 18 AND Y = 10 else
"1111111111111" when X = 19 AND Y = 10 else
"1111111111111" when X = 20 AND Y = 10 else
"1111111111111" when X = 21 AND Y = 10 else
"1111111111111" when X = 22 AND Y = 10 else
"1111111111111" when X = 23 AND Y = 10 else
"1111111111111" when X = 24 AND Y = 10 else
"1111111111111" when X = 25 AND Y = 10 else
"1111111111111" when X = 26 AND Y = 10 else
"1111111111111" when X = 27 AND Y = 10 else
"1111111111111" when X = 28 AND Y = 10 else
"1111111111111" when X = 29 AND Y = 10 else
"1111111111111" when X = 30 AND Y = 10 else
"1111111111111" when X = 31 AND Y = 10 else
"1111111111111" when X = 32 AND Y = 10 else
"1111111111111" when X = 33 AND Y = 10 else
"1111111111111" when X = 34 AND Y = 10 else
"1111111111111" when X = 35 AND Y = 10 else
"1111111111111" when X = 36 AND Y = 10 else
"1111111111111" when X = 37 AND Y = 10 else
"1111111111111" when X = 38 AND Y = 10 else
"1111111111111" when X = 39 AND Y = 10 else
"1111111111111" when X = 40 AND Y = 10 else
"1111111111111" when X = 41 AND Y = 10 else
"1111111111111" when X = 42 AND Y = 10 else
"1111111111111" when X = 43 AND Y = 10 else
"1111111111111" when X = 44 AND Y = 10 else
"1111111111111" when X = 45 AND Y = 10 else
"1111111111111" when X = 46 AND Y = 10 else
"1111111111111" when X = 47 AND Y = 10 else
"1111111111111" when X = 48 AND Y = 10 else
"1111111111111" when X = 49 AND Y = 10 else
"1111111111111" when X = 50 AND Y = 10 else
"1111111111111" when X = 51 AND Y = 10 else
"1111111111111" when X = 52 AND Y = 10 else
"1111111111111" when X = 53 AND Y = 10 else
"1111111111111" when X = 54 AND Y = 10 else
"1111111111111" when X = 55 AND Y = 10 else
"1111111111111" when X = 56 AND Y = 10 else
"1111111111111" when X = 57 AND Y = 10 else
"1111111111111" when X = 58 AND Y = 10 else
"1111111111111" when X = 59 AND Y = 10 else
"1111111111111" when X = 60 AND Y = 10 else
"1101111011111" when X = 61 AND Y = 10 else
"1101110111111" when X = 62 AND Y = 10 else
"1101110111111" when X = 63 AND Y = 10 else
"1010101011001" when X = 64 AND Y = 10 else
"0000000000000" when X = 65 AND Y = 10 else
"0000000000000" when X = 66 AND Y = 10 else
"0000000000000" when X = 67 AND Y = 10 else
"0000000000000" when X = 68 AND Y = 10 else
"0000000000000" when X = 69 AND Y = 10 else
"0000000000000" when X = 70 AND Y = 10 else
"0000000000000" when X = 71 AND Y = 10 else
"0000000000000" when X = 72 AND Y = 10 else
"0000000000000" when X = 73 AND Y = 10 else
"0000000000000" when X = 74 AND Y = 10 else
"0000000000000" when X = 0 AND Y = 11 else
"0000000000000" when X = 1 AND Y = 11 else
"0000000000000" when X = 2 AND Y = 11 else
"0000000000000" when X = 3 AND Y = 11 else
"0000000000000" when X = 4 AND Y = 11 else
"0000000000000" when X = 5 AND Y = 11 else
"0000000000000" when X = 6 AND Y = 11 else
"0001000100101" when X = 7 AND Y = 11 else
"0101011010011" when X = 8 AND Y = 11 else
"0101011010101" when X = 9 AND Y = 11 else
"1001100111001" when X = 10 AND Y = 11 else
"1100110011101" when X = 11 AND Y = 11 else
"1101110111111" when X = 12 AND Y = 11 else
"1101110111111" when X = 13 AND Y = 11 else
"1110111011111" when X = 14 AND Y = 11 else
"1110111011111" when X = 15 AND Y = 11 else
"1111111111111" when X = 16 AND Y = 11 else
"1111111111111" when X = 17 AND Y = 11 else
"1111111111111" when X = 18 AND Y = 11 else
"1111111111111" when X = 19 AND Y = 11 else
"1111111111111" when X = 20 AND Y = 11 else
"1111111111111" when X = 21 AND Y = 11 else
"1111111111111" when X = 22 AND Y = 11 else
"1111111111111" when X = 23 AND Y = 11 else
"1111111111111" when X = 24 AND Y = 11 else
"1111111111111" when X = 25 AND Y = 11 else
"1111111111111" when X = 26 AND Y = 11 else
"1111111111111" when X = 27 AND Y = 11 else
"1111111111111" when X = 28 AND Y = 11 else
"1111111111111" when X = 29 AND Y = 11 else
"1111111111111" when X = 30 AND Y = 11 else
"1111111111111" when X = 31 AND Y = 11 else
"1111111111111" when X = 32 AND Y = 11 else
"1111111111111" when X = 33 AND Y = 11 else
"1111111111111" when X = 34 AND Y = 11 else
"1111111111111" when X = 35 AND Y = 11 else
"1111111111111" when X = 36 AND Y = 11 else
"1111111111111" when X = 37 AND Y = 11 else
"1111111111111" when X = 38 AND Y = 11 else
"1111111111111" when X = 39 AND Y = 11 else
"1111111111111" when X = 40 AND Y = 11 else
"1111111111111" when X = 41 AND Y = 11 else
"1111111111111" when X = 42 AND Y = 11 else
"1111111111111" when X = 43 AND Y = 11 else
"1111111111111" when X = 44 AND Y = 11 else
"1111111111111" when X = 45 AND Y = 11 else
"1111111111111" when X = 46 AND Y = 11 else
"1111111111111" when X = 47 AND Y = 11 else
"1111111111111" when X = 48 AND Y = 11 else
"1111111111111" when X = 49 AND Y = 11 else
"1111111111111" when X = 50 AND Y = 11 else
"1111111111111" when X = 51 AND Y = 11 else
"1111111111111" when X = 52 AND Y = 11 else
"1111111111111" when X = 53 AND Y = 11 else
"1111111111111" when X = 54 AND Y = 11 else
"1111111111111" when X = 55 AND Y = 11 else
"1111111111111" when X = 56 AND Y = 11 else
"1111111111111" when X = 57 AND Y = 11 else
"1111111111111" when X = 58 AND Y = 11 else
"1111111111111" when X = 59 AND Y = 11 else
"1111111111111" when X = 60 AND Y = 11 else
"1101111011111" when X = 61 AND Y = 11 else
"1101110111111" when X = 62 AND Y = 11 else
"1101110111111" when X = 63 AND Y = 11 else
"1010101011001" when X = 64 AND Y = 11 else
"0000000000000" when X = 65 AND Y = 11 else
"0000000000000" when X = 66 AND Y = 11 else
"0000000000000" when X = 67 AND Y = 11 else
"0000000000000" when X = 68 AND Y = 11 else
"0000000000000" when X = 69 AND Y = 11 else
"0000000000000" when X = 70 AND Y = 11 else
"0000000000000" when X = 71 AND Y = 11 else
"0000000000000" when X = 72 AND Y = 11 else
"0000000000000" when X = 73 AND Y = 11 else
"0000000000000" when X = 74 AND Y = 11 else
"0000000000000" when X = 0 AND Y = 12 else
"0000000000000" when X = 1 AND Y = 12 else
"0000000000000" when X = 2 AND Y = 12 else
"0000000000000" when X = 3 AND Y = 12 else
"0000000000000" when X = 4 AND Y = 12 else
"0000000000000" when X = 5 AND Y = 12 else
"0001001000111" when X = 6 AND Y = 12 else
"0101011010011" when X = 7 AND Y = 12 else
"0111100011011" when X = 8 AND Y = 12 else
"1001101011101" when X = 9 AND Y = 12 else
"1100110011101" when X = 10 AND Y = 12 else
"1101110111111" when X = 11 AND Y = 12 else
"1101110111111" when X = 12 AND Y = 12 else
"1101110111111" when X = 13 AND Y = 12 else
"1101110111111" when X = 14 AND Y = 12 else
"1101110111111" when X = 15 AND Y = 12 else
"1110111011111" when X = 16 AND Y = 12 else
"1110111111111" when X = 17 AND Y = 12 else
"1110111111111" when X = 18 AND Y = 12 else
"1110111111111" when X = 19 AND Y = 12 else
"1110111111111" when X = 20 AND Y = 12 else
"1111111111111" when X = 21 AND Y = 12 else
"1111111111111" when X = 22 AND Y = 12 else
"1111111111111" when X = 23 AND Y = 12 else
"1111111111111" when X = 24 AND Y = 12 else
"1111111111111" when X = 25 AND Y = 12 else
"1111111111111" when X = 26 AND Y = 12 else
"1111111111111" when X = 27 AND Y = 12 else
"1111111111111" when X = 28 AND Y = 12 else
"1111111111111" when X = 29 AND Y = 12 else
"1111111111111" when X = 30 AND Y = 12 else
"1111111111111" when X = 31 AND Y = 12 else
"1111111111111" when X = 32 AND Y = 12 else
"1111111111111" when X = 33 AND Y = 12 else
"1111111111111" when X = 34 AND Y = 12 else
"1111111111111" when X = 35 AND Y = 12 else
"1111111111111" when X = 36 AND Y = 12 else
"1111111111111" when X = 37 AND Y = 12 else
"1111111111111" when X = 38 AND Y = 12 else
"1111111111111" when X = 39 AND Y = 12 else
"1111111111111" when X = 40 AND Y = 12 else
"1111111111111" when X = 41 AND Y = 12 else
"1111111111111" when X = 42 AND Y = 12 else
"1111111111111" when X = 43 AND Y = 12 else
"1111111111111" when X = 44 AND Y = 12 else
"1111111111111" when X = 45 AND Y = 12 else
"1111111111111" when X = 46 AND Y = 12 else
"1111111111111" when X = 47 AND Y = 12 else
"1111111111111" when X = 48 AND Y = 12 else
"1111111111111" when X = 49 AND Y = 12 else
"1111111111111" when X = 50 AND Y = 12 else
"1111111111111" when X = 51 AND Y = 12 else
"1111111111111" when X = 52 AND Y = 12 else
"1111111111111" when X = 53 AND Y = 12 else
"1111111111111" when X = 54 AND Y = 12 else
"1111111111111" when X = 55 AND Y = 12 else
"1111111111111" when X = 56 AND Y = 12 else
"1111111111111" when X = 57 AND Y = 12 else
"1111111111111" when X = 58 AND Y = 12 else
"1111111111111" when X = 59 AND Y = 12 else
"1111111111111" when X = 60 AND Y = 12 else
"1101111011111" when X = 61 AND Y = 12 else
"1101110111111" when X = 62 AND Y = 12 else
"1101110111111" when X = 63 AND Y = 12 else
"1010101011001" when X = 64 AND Y = 12 else
"0000000000000" when X = 65 AND Y = 12 else
"0000000000000" when X = 66 AND Y = 12 else
"0000000000000" when X = 67 AND Y = 12 else
"0000000000000" when X = 68 AND Y = 12 else
"0000000000000" when X = 69 AND Y = 12 else
"0000000000000" when X = 70 AND Y = 12 else
"0000000000000" when X = 71 AND Y = 12 else
"0000000000000" when X = 72 AND Y = 12 else
"0000000000000" when X = 73 AND Y = 12 else
"0000000000000" when X = 74 AND Y = 12 else
"0000000000000" when X = 0 AND Y = 13 else
"0000000000000" when X = 1 AND Y = 13 else
"0000000000000" when X = 2 AND Y = 13 else
"0000000000000" when X = 3 AND Y = 13 else
"0000000000000" when X = 4 AND Y = 13 else
"0010001000111" when X = 5 AND Y = 13 else
"0101010110001" when X = 6 AND Y = 13 else
"1000100111011" when X = 7 AND Y = 13 else
"1001101011101" when X = 8 AND Y = 13 else
"1100110011101" when X = 9 AND Y = 13 else
"1101110111111" when X = 10 AND Y = 13 else
"1101110111111" when X = 11 AND Y = 13 else
"1101110111111" when X = 12 AND Y = 13 else
"1101110111111" when X = 13 AND Y = 13 else
"1101110111111" when X = 14 AND Y = 13 else
"1101110111111" when X = 15 AND Y = 13 else
"1101110111111" when X = 16 AND Y = 13 else
"1101110111111" when X = 17 AND Y = 13 else
"1101110111111" when X = 18 AND Y = 13 else
"1101110111111" when X = 19 AND Y = 13 else
"1101110111111" when X = 20 AND Y = 13 else
"1101110111111" when X = 21 AND Y = 13 else
"1111111111111" when X = 22 AND Y = 13 else
"1111111111111" when X = 23 AND Y = 13 else
"1111111111111" when X = 24 AND Y = 13 else
"1111111111111" when X = 25 AND Y = 13 else
"1111111111111" when X = 26 AND Y = 13 else
"1111111111111" when X = 27 AND Y = 13 else
"1111111111111" when X = 28 AND Y = 13 else
"1111111111111" when X = 29 AND Y = 13 else
"1111111111111" when X = 30 AND Y = 13 else
"1111111111111" when X = 31 AND Y = 13 else
"1111111111111" when X = 32 AND Y = 13 else
"1111111111111" when X = 33 AND Y = 13 else
"1111111111111" when X = 34 AND Y = 13 else
"1111111111111" when X = 35 AND Y = 13 else
"1111111111111" when X = 36 AND Y = 13 else
"1111111111111" when X = 37 AND Y = 13 else
"1111111111111" when X = 38 AND Y = 13 else
"1111111111111" when X = 39 AND Y = 13 else
"1111111111111" when X = 40 AND Y = 13 else
"1111111111111" when X = 41 AND Y = 13 else
"1111111111111" when X = 42 AND Y = 13 else
"1111111111111" when X = 43 AND Y = 13 else
"1111111111111" when X = 44 AND Y = 13 else
"1111111111111" when X = 45 AND Y = 13 else
"1111111111111" when X = 46 AND Y = 13 else
"1111111111111" when X = 47 AND Y = 13 else
"1111111111111" when X = 48 AND Y = 13 else
"1111111111111" when X = 49 AND Y = 13 else
"1111111111111" when X = 50 AND Y = 13 else
"1111111111111" when X = 51 AND Y = 13 else
"1111111111111" when X = 52 AND Y = 13 else
"1111111111111" when X = 53 AND Y = 13 else
"1111111111111" when X = 54 AND Y = 13 else
"1111111111111" when X = 55 AND Y = 13 else
"1111111111111" when X = 56 AND Y = 13 else
"1111111111111" when X = 57 AND Y = 13 else
"1111111111111" when X = 58 AND Y = 13 else
"1111111111111" when X = 59 AND Y = 13 else
"1111111111111" when X = 60 AND Y = 13 else
"1101111011111" when X = 61 AND Y = 13 else
"1101110111111" when X = 62 AND Y = 13 else
"1101110111111" when X = 63 AND Y = 13 else
"1010101011001" when X = 64 AND Y = 13 else
"0000000000000" when X = 65 AND Y = 13 else
"0000000000000" when X = 66 AND Y = 13 else
"0000000000000" when X = 67 AND Y = 13 else
"0000000000000" when X = 68 AND Y = 13 else
"0000000000000" when X = 69 AND Y = 13 else
"0000000000000" when X = 70 AND Y = 13 else
"0000000000000" when X = 71 AND Y = 13 else
"0000000000000" when X = 72 AND Y = 13 else
"0000000000000" when X = 73 AND Y = 13 else
"0000000000000" when X = 74 AND Y = 13 else
"0000000000000" when X = 0 AND Y = 14 else
"0000000000000" when X = 1 AND Y = 14 else
"0000000000000" when X = 2 AND Y = 14 else
"0000000000000" when X = 3 AND Y = 14 else
"0010001000111" when X = 4 AND Y = 14 else
"0101010110001" when X = 5 AND Y = 14 else
"0111100111011" when X = 6 AND Y = 14 else
"1000100111011" when X = 7 AND Y = 14 else
"1100110011101" when X = 8 AND Y = 14 else
"1101110111111" when X = 9 AND Y = 14 else
"1101110111111" when X = 10 AND Y = 14 else
"1101110111111" when X = 11 AND Y = 14 else
"1101110111111" when X = 12 AND Y = 14 else
"1101110111111" when X = 13 AND Y = 14 else
"1101110111111" when X = 14 AND Y = 14 else
"1101110111111" when X = 15 AND Y = 14 else
"1101110111111" when X = 16 AND Y = 14 else
"1101110111111" when X = 17 AND Y = 14 else
"1101110111111" when X = 18 AND Y = 14 else
"1101110111111" when X = 19 AND Y = 14 else
"1101110111111" when X = 20 AND Y = 14 else
"1101110111111" when X = 21 AND Y = 14 else
"1101110111111" when X = 22 AND Y = 14 else
"1111111111111" when X = 23 AND Y = 14 else
"1111111111111" when X = 24 AND Y = 14 else
"1111111111111" when X = 25 AND Y = 14 else
"1111111111111" when X = 26 AND Y = 14 else
"1111111111111" when X = 27 AND Y = 14 else
"1111111111111" when X = 28 AND Y = 14 else
"1111111111111" when X = 29 AND Y = 14 else
"1111111111111" when X = 30 AND Y = 14 else
"1111111111111" when X = 31 AND Y = 14 else
"1111111111111" when X = 32 AND Y = 14 else
"1111111111111" when X = 33 AND Y = 14 else
"1111111111111" when X = 34 AND Y = 14 else
"1111111111111" when X = 35 AND Y = 14 else
"1111111111111" when X = 36 AND Y = 14 else
"1111111111111" when X = 37 AND Y = 14 else
"1111111111111" when X = 38 AND Y = 14 else
"1111111111111" when X = 39 AND Y = 14 else
"1111111111111" when X = 40 AND Y = 14 else
"1111111111111" when X = 41 AND Y = 14 else
"1111111111111" when X = 42 AND Y = 14 else
"1111111111111" when X = 43 AND Y = 14 else
"1111111111111" when X = 44 AND Y = 14 else
"1111111111111" when X = 45 AND Y = 14 else
"1111111111111" when X = 46 AND Y = 14 else
"1111111111111" when X = 47 AND Y = 14 else
"1111111111111" when X = 48 AND Y = 14 else
"1111111111111" when X = 49 AND Y = 14 else
"1111111111111" when X = 50 AND Y = 14 else
"1111111111111" when X = 51 AND Y = 14 else
"1111111111111" when X = 52 AND Y = 14 else
"1111111111111" when X = 53 AND Y = 14 else
"1111111111111" when X = 54 AND Y = 14 else
"1111111111111" when X = 55 AND Y = 14 else
"1111111111111" when X = 56 AND Y = 14 else
"1111111111111" when X = 57 AND Y = 14 else
"1111111111111" when X = 58 AND Y = 14 else
"1111111111111" when X = 59 AND Y = 14 else
"1111111111111" when X = 60 AND Y = 14 else
"1101111011111" when X = 61 AND Y = 14 else
"1101110111111" when X = 62 AND Y = 14 else
"1101110111111" when X = 63 AND Y = 14 else
"1010101011001" when X = 64 AND Y = 14 else
"0000000000000" when X = 65 AND Y = 14 else
"0000000000000" when X = 66 AND Y = 14 else
"0000000000000" when X = 67 AND Y = 14 else
"0000000000000" when X = 68 AND Y = 14 else
"0000000000000" when X = 69 AND Y = 14 else
"0000000000000" when X = 70 AND Y = 14 else
"0000000000000" when X = 71 AND Y = 14 else
"0000000000000" when X = 72 AND Y = 14 else
"0000000000000" when X = 73 AND Y = 14 else
"0000000000000" when X = 74 AND Y = 14 else
"0000000000000" when X = 0 AND Y = 15 else
"0000000000000" when X = 1 AND Y = 15 else
"0001001000111" when X = 2 AND Y = 15 else
"0010001001001" when X = 3 AND Y = 15 else
"0101011010011" when X = 4 AND Y = 15 else
"0111100011011" when X = 5 AND Y = 15 else
"1000100111011" when X = 6 AND Y = 15 else
"1000100111011" when X = 7 AND Y = 15 else
"1100110111101" when X = 8 AND Y = 15 else
"1101110111111" when X = 9 AND Y = 15 else
"1101110111111" when X = 10 AND Y = 15 else
"1101110111111" when X = 11 AND Y = 15 else
"1101110111111" when X = 12 AND Y = 15 else
"1101110111111" when X = 13 AND Y = 15 else
"1101110111111" when X = 14 AND Y = 15 else
"1101110111111" when X = 15 AND Y = 15 else
"1101110111111" when X = 16 AND Y = 15 else
"1101110111111" when X = 17 AND Y = 15 else
"1101110111111" when X = 18 AND Y = 15 else
"1101110111111" when X = 19 AND Y = 15 else
"1101110111111" when X = 20 AND Y = 15 else
"1101110111111" when X = 21 AND Y = 15 else
"1101110111111" when X = 22 AND Y = 15 else
"1101110111111" when X = 23 AND Y = 15 else
"1111111111111" when X = 24 AND Y = 15 else
"1111111111111" when X = 25 AND Y = 15 else
"1111111111111" when X = 26 AND Y = 15 else
"1111111111111" when X = 27 AND Y = 15 else
"1111111111111" when X = 28 AND Y = 15 else
"1111111111111" when X = 29 AND Y = 15 else
"1111111111111" when X = 30 AND Y = 15 else
"1111111111111" when X = 31 AND Y = 15 else
"1111111111111" when X = 32 AND Y = 15 else
"1111111111111" when X = 33 AND Y = 15 else
"1111111111111" when X = 34 AND Y = 15 else
"1111111111111" when X = 35 AND Y = 15 else
"1111111111111" when X = 36 AND Y = 15 else
"1111111111111" when X = 37 AND Y = 15 else
"1111111111111" when X = 38 AND Y = 15 else
"1111111111111" when X = 39 AND Y = 15 else
"1111111111111" when X = 40 AND Y = 15 else
"1111111111111" when X = 41 AND Y = 15 else
"1111111111111" when X = 42 AND Y = 15 else
"1111111111111" when X = 43 AND Y = 15 else
"1111111111111" when X = 44 AND Y = 15 else
"1111111111111" when X = 45 AND Y = 15 else
"1111111111111" when X = 46 AND Y = 15 else
"1111111111111" when X = 47 AND Y = 15 else
"1111111111111" when X = 48 AND Y = 15 else
"1111111111111" when X = 49 AND Y = 15 else
"1111111111111" when X = 50 AND Y = 15 else
"1111111111111" when X = 51 AND Y = 15 else
"1111111111111" when X = 52 AND Y = 15 else
"1111111111111" when X = 53 AND Y = 15 else
"1111111111111" when X = 54 AND Y = 15 else
"1111111111111" when X = 55 AND Y = 15 else
"1111111111111" when X = 56 AND Y = 15 else
"1111111111111" when X = 57 AND Y = 15 else
"1111111111111" when X = 58 AND Y = 15 else
"1111111111111" when X = 59 AND Y = 15 else
"1111111111111" when X = 60 AND Y = 15 else
"1101111011111" when X = 61 AND Y = 15 else
"1101110111111" when X = 62 AND Y = 15 else
"1101110111111" when X = 63 AND Y = 15 else
"1010101011001" when X = 64 AND Y = 15 else
"0000000000000" when X = 65 AND Y = 15 else
"0000000000000" when X = 66 AND Y = 15 else
"0000000000000" when X = 67 AND Y = 15 else
"0000000000000" when X = 68 AND Y = 15 else
"0000000000000" when X = 69 AND Y = 15 else
"0000000000000" when X = 70 AND Y = 15 else
"0000000000000" when X = 71 AND Y = 15 else
"0000000000000" when X = 72 AND Y = 15 else
"0000000000000" when X = 73 AND Y = 15 else
"0000000000000" when X = 74 AND Y = 15 else
"0000000000000" when X = 0 AND Y = 16 else
"0001000100101" when X = 1 AND Y = 16 else
"0110011110101" when X = 2 AND Y = 16 else
"0111100011001" when X = 3 AND Y = 16 else
"0111100011011" when X = 4 AND Y = 16 else
"1000100111011" when X = 5 AND Y = 16 else
"1000100111011" when X = 6 AND Y = 16 else
"1100110011101" when X = 7 AND Y = 16 else
"1101110111111" when X = 8 AND Y = 16 else
"1101110111111" when X = 9 AND Y = 16 else
"1101110111111" when X = 10 AND Y = 16 else
"1101110111111" when X = 11 AND Y = 16 else
"1101110111111" when X = 12 AND Y = 16 else
"1101110111111" when X = 13 AND Y = 16 else
"1101110111111" when X = 14 AND Y = 16 else
"1101110111111" when X = 15 AND Y = 16 else
"1101110111111" when X = 16 AND Y = 16 else
"1101110111111" when X = 17 AND Y = 16 else
"1101110111111" when X = 18 AND Y = 16 else
"1101110111111" when X = 19 AND Y = 16 else
"1101110111111" when X = 20 AND Y = 16 else
"1101110111111" when X = 21 AND Y = 16 else
"1101110111111" when X = 22 AND Y = 16 else
"1101110111111" when X = 23 AND Y = 16 else
"1111111111111" when X = 24 AND Y = 16 else
"1111111111111" when X = 25 AND Y = 16 else
"1111111111111" when X = 26 AND Y = 16 else
"1111111111111" when X = 27 AND Y = 16 else
"1111111111111" when X = 28 AND Y = 16 else
"1111111111111" when X = 29 AND Y = 16 else
"1111111111111" when X = 30 AND Y = 16 else
"1111111111111" when X = 31 AND Y = 16 else
"1111111111111" when X = 32 AND Y = 16 else
"1111111111111" when X = 33 AND Y = 16 else
"1111111111111" when X = 34 AND Y = 16 else
"1111111111111" when X = 35 AND Y = 16 else
"1111111111111" when X = 36 AND Y = 16 else
"1111111111111" when X = 37 AND Y = 16 else
"1111111111111" when X = 38 AND Y = 16 else
"1111111111111" when X = 39 AND Y = 16 else
"1111111111111" when X = 40 AND Y = 16 else
"1111111111111" when X = 41 AND Y = 16 else
"1111111111111" when X = 42 AND Y = 16 else
"1111111111111" when X = 43 AND Y = 16 else
"1111111111111" when X = 44 AND Y = 16 else
"1111111111111" when X = 45 AND Y = 16 else
"1111111111111" when X = 46 AND Y = 16 else
"1111111111111" when X = 47 AND Y = 16 else
"1111111111111" when X = 48 AND Y = 16 else
"1111111111111" when X = 49 AND Y = 16 else
"1111111111111" when X = 50 AND Y = 16 else
"1111111111111" when X = 51 AND Y = 16 else
"1111111111111" when X = 52 AND Y = 16 else
"1111111111111" when X = 53 AND Y = 16 else
"1111111111111" when X = 54 AND Y = 16 else
"1111111111111" when X = 55 AND Y = 16 else
"1111111111111" when X = 56 AND Y = 16 else
"1111111111111" when X = 57 AND Y = 16 else
"1111111111111" when X = 58 AND Y = 16 else
"1111111111111" when X = 59 AND Y = 16 else
"1111111111111" when X = 60 AND Y = 16 else
"1101111011111" when X = 61 AND Y = 16 else
"1101110111111" when X = 62 AND Y = 16 else
"1101110111101" when X = 63 AND Y = 16 else
"1010101010111" when X = 64 AND Y = 16 else
"0000000000000" when X = 65 AND Y = 16 else
"0000000000000" when X = 66 AND Y = 16 else
"0000000000000" when X = 67 AND Y = 16 else
"0000000000000" when X = 68 AND Y = 16 else
"0000000000000" when X = 69 AND Y = 16 else
"0000000000000" when X = 70 AND Y = 16 else
"0000000000000" when X = 71 AND Y = 16 else
"0000000000000" when X = 72 AND Y = 16 else
"0000000000000" when X = 73 AND Y = 16 else
"0000000000000" when X = 74 AND Y = 16 else
"0001000100101" when X = 0 AND Y = 17 else
"0110011110101" when X = 1 AND Y = 17 else
"0111100011011" when X = 2 AND Y = 17 else
"1000100111011" when X = 3 AND Y = 17 else
"1000100111011" when X = 4 AND Y = 17 else
"1000100111011" when X = 5 AND Y = 17 else
"1001100111011" when X = 6 AND Y = 17 else
"1101110111101" when X = 7 AND Y = 17 else
"1101110111111" when X = 8 AND Y = 17 else
"1101110111111" when X = 9 AND Y = 17 else
"1101110111111" when X = 10 AND Y = 17 else
"1101110111111" when X = 11 AND Y = 17 else
"1101110111111" when X = 12 AND Y = 17 else
"1101110111111" when X = 13 AND Y = 17 else
"1101110111111" when X = 14 AND Y = 17 else
"1101110111111" when X = 15 AND Y = 17 else
"1101110111111" when X = 16 AND Y = 17 else
"1101110111111" when X = 17 AND Y = 17 else
"1101110111111" when X = 18 AND Y = 17 else
"1101110111111" when X = 19 AND Y = 17 else
"1101110111111" when X = 20 AND Y = 17 else
"1101110111111" when X = 21 AND Y = 17 else
"1101110111111" when X = 22 AND Y = 17 else
"1101110111111" when X = 23 AND Y = 17 else
"1101111011111" when X = 24 AND Y = 17 else
"1111111111111" when X = 25 AND Y = 17 else
"1111111111111" when X = 26 AND Y = 17 else
"1111111111111" when X = 27 AND Y = 17 else
"1111111111111" when X = 28 AND Y = 17 else
"1111111111111" when X = 29 AND Y = 17 else
"1111111111111" when X = 30 AND Y = 17 else
"1111111111111" when X = 31 AND Y = 17 else
"1111111111111" when X = 32 AND Y = 17 else
"1111111111111" when X = 33 AND Y = 17 else
"1111111111111" when X = 34 AND Y = 17 else
"1111111111111" when X = 35 AND Y = 17 else
"1111111111111" when X = 36 AND Y = 17 else
"1111111111111" when X = 37 AND Y = 17 else
"1111111111111" when X = 38 AND Y = 17 else
"1111111111111" when X = 39 AND Y = 17 else
"1111111111111" when X = 40 AND Y = 17 else
"1111111111111" when X = 41 AND Y = 17 else
"1111111111111" when X = 42 AND Y = 17 else
"1111111111111" when X = 43 AND Y = 17 else
"1111111111111" when X = 44 AND Y = 17 else
"1111111111111" when X = 45 AND Y = 17 else
"1111111111111" when X = 46 AND Y = 17 else
"1111111111111" when X = 47 AND Y = 17 else
"1111111111111" when X = 48 AND Y = 17 else
"1111111111111" when X = 49 AND Y = 17 else
"1111111111111" when X = 50 AND Y = 17 else
"1111111111111" when X = 51 AND Y = 17 else
"1111111111111" when X = 52 AND Y = 17 else
"1111111111111" when X = 53 AND Y = 17 else
"1111111111111" when X = 54 AND Y = 17 else
"1111111111111" when X = 55 AND Y = 17 else
"1111111111111" when X = 56 AND Y = 17 else
"1111111111111" when X = 57 AND Y = 17 else
"1111111111111" when X = 58 AND Y = 17 else
"1111111111111" when X = 59 AND Y = 17 else
"1111111111111" when X = 60 AND Y = 17 else
"1101111011111" when X = 61 AND Y = 17 else
"1101110111111" when X = 62 AND Y = 17 else
"1010101011001" when X = 63 AND Y = 17 else
"0101010101101" when X = 64 AND Y = 17 else
"0000000000000" when X = 65 AND Y = 17 else
"0000000000000" when X = 66 AND Y = 17 else
"0000000000000" when X = 67 AND Y = 17 else
"0000000000000" when X = 68 AND Y = 17 else
"0000000000000" when X = 69 AND Y = 17 else
"0000000000000" when X = 70 AND Y = 17 else
"0000000000000" when X = 71 AND Y = 17 else
"0000000000000" when X = 72 AND Y = 17 else
"0000000000000" when X = 73 AND Y = 17 else
"0000000000000" when X = 74 AND Y = 17 else
"0110011110111" when X = 0 AND Y = 18 else
"0111100011011" when X = 1 AND Y = 18 else
"1000100111011" when X = 2 AND Y = 18 else
"1000100111011" when X = 3 AND Y = 18 else
"1000100111011" when X = 4 AND Y = 18 else
"1000100111011" when X = 5 AND Y = 18 else
"1000100111011" when X = 6 AND Y = 18 else
"1100110111101" when X = 7 AND Y = 18 else
"1101110111111" when X = 8 AND Y = 18 else
"1101110111111" when X = 9 AND Y = 18 else
"1101110111111" when X = 10 AND Y = 18 else
"1101110111111" when X = 11 AND Y = 18 else
"1101110111111" when X = 12 AND Y = 18 else
"1101110111111" when X = 13 AND Y = 18 else
"1101110111111" when X = 14 AND Y = 18 else
"1101110111111" when X = 15 AND Y = 18 else
"1101110111111" when X = 16 AND Y = 18 else
"1101110111111" when X = 17 AND Y = 18 else
"1101110111111" when X = 18 AND Y = 18 else
"1101110111111" when X = 19 AND Y = 18 else
"1101110111111" when X = 20 AND Y = 18 else
"1101110111111" when X = 21 AND Y = 18 else
"1101110111111" when X = 22 AND Y = 18 else
"1101110111111" when X = 23 AND Y = 18 else
"1110111011111" when X = 24 AND Y = 18 else
"1111111111111" when X = 25 AND Y = 18 else
"1111111111111" when X = 26 AND Y = 18 else
"1111111111111" when X = 27 AND Y = 18 else
"1111111111111" when X = 28 AND Y = 18 else
"1111111111111" when X = 29 AND Y = 18 else
"1111111111111" when X = 30 AND Y = 18 else
"1111111111111" when X = 31 AND Y = 18 else
"1111111111111" when X = 32 AND Y = 18 else
"1111111111111" when X = 33 AND Y = 18 else
"1111111111111" when X = 34 AND Y = 18 else
"1111111111111" when X = 35 AND Y = 18 else
"1111111111111" when X = 36 AND Y = 18 else
"1111111111111" when X = 37 AND Y = 18 else
"1111111111111" when X = 38 AND Y = 18 else
"1111111111111" when X = 39 AND Y = 18 else
"1111111111111" when X = 40 AND Y = 18 else
"1111111111111" when X = 41 AND Y = 18 else
"1111111111111" when X = 42 AND Y = 18 else
"1111111111111" when X = 43 AND Y = 18 else
"1111111111111" when X = 44 AND Y = 18 else
"1111111111111" when X = 45 AND Y = 18 else
"1111111111111" when X = 46 AND Y = 18 else
"1111111111111" when X = 47 AND Y = 18 else
"1111111111111" when X = 48 AND Y = 18 else
"1111111111111" when X = 49 AND Y = 18 else
"1111111111111" when X = 50 AND Y = 18 else
"1111111111111" when X = 51 AND Y = 18 else
"1111111111111" when X = 52 AND Y = 18 else
"1111111111111" when X = 53 AND Y = 18 else
"1111111111111" when X = 54 AND Y = 18 else
"1111111111111" when X = 55 AND Y = 18 else
"1111111111111" when X = 56 AND Y = 18 else
"1111111111111" when X = 57 AND Y = 18 else
"1111111111111" when X = 58 AND Y = 18 else
"1111111111111" when X = 59 AND Y = 18 else
"1111111111111" when X = 60 AND Y = 18 else
"1111111111111" when X = 61 AND Y = 18 else
"1101111011111" when X = 62 AND Y = 18 else
"1011110011011" when X = 63 AND Y = 18 else
"1010101011001" when X = 64 AND Y = 18 else
"1001100110101" when X = 65 AND Y = 18 else
"0000000000000" when X = 66 AND Y = 18 else
"0000000000000" when X = 67 AND Y = 18 else
"0000000000000" when X = 68 AND Y = 18 else
"0000000000000" when X = 69 AND Y = 18 else
"0000000000000" when X = 70 AND Y = 18 else
"0000000000000" when X = 71 AND Y = 18 else
"0000000000000" when X = 72 AND Y = 18 else
"0000000000000" when X = 73 AND Y = 18 else
"0000000000000" when X = 74 AND Y = 18 else
"1000100111011" when X = 0 AND Y = 19 else
"1000100111011" when X = 1 AND Y = 19 else
"1000100111011" when X = 2 AND Y = 19 else
"1000100111011" when X = 3 AND Y = 19 else
"1000100111011" when X = 4 AND Y = 19 else
"1000100111011" when X = 5 AND Y = 19 else
"1011101111101" when X = 6 AND Y = 19 else
"1101110111111" when X = 7 AND Y = 19 else
"1101110111111" when X = 8 AND Y = 19 else
"1101110111111" when X = 9 AND Y = 19 else
"1101110111111" when X = 10 AND Y = 19 else
"1101110111111" when X = 11 AND Y = 19 else
"1101110111111" when X = 12 AND Y = 19 else
"1101110111111" when X = 13 AND Y = 19 else
"1101110111111" when X = 14 AND Y = 19 else
"1101110111111" when X = 15 AND Y = 19 else
"1101110111111" when X = 16 AND Y = 19 else
"1101110111111" when X = 17 AND Y = 19 else
"1101110111111" when X = 18 AND Y = 19 else
"1101110111111" when X = 19 AND Y = 19 else
"1101110111111" when X = 20 AND Y = 19 else
"1101110111111" when X = 21 AND Y = 19 else
"1101110111111" when X = 22 AND Y = 19 else
"1110111011111" when X = 23 AND Y = 19 else
"1111111111111" when X = 24 AND Y = 19 else
"1111111111111" when X = 25 AND Y = 19 else
"1111111111111" when X = 26 AND Y = 19 else
"1111111111111" when X = 27 AND Y = 19 else
"1111111111111" when X = 28 AND Y = 19 else
"1111111111111" when X = 29 AND Y = 19 else
"1111111111111" when X = 30 AND Y = 19 else
"1111111111111" when X = 31 AND Y = 19 else
"1111111111111" when X = 32 AND Y = 19 else
"1111111111111" when X = 33 AND Y = 19 else
"1111111111111" when X = 34 AND Y = 19 else
"1111111111111" when X = 35 AND Y = 19 else
"1111111111111" when X = 36 AND Y = 19 else
"1111111111111" when X = 37 AND Y = 19 else
"1111111111111" when X = 38 AND Y = 19 else
"1111111111111" when X = 39 AND Y = 19 else
"1111111111111" when X = 40 AND Y = 19 else
"1111111111111" when X = 41 AND Y = 19 else
"1111111111111" when X = 42 AND Y = 19 else
"1111111111111" when X = 43 AND Y = 19 else
"1111111111111" when X = 44 AND Y = 19 else
"1111111111111" when X = 45 AND Y = 19 else
"1111111111111" when X = 46 AND Y = 19 else
"1111111111111" when X = 47 AND Y = 19 else
"1111111111111" when X = 48 AND Y = 19 else
"1111111111111" when X = 49 AND Y = 19 else
"1111111111111" when X = 50 AND Y = 19 else
"1111111111111" when X = 51 AND Y = 19 else
"1111111111111" when X = 52 AND Y = 19 else
"1111111111111" when X = 53 AND Y = 19 else
"1111111111111" when X = 54 AND Y = 19 else
"1111111111111" when X = 55 AND Y = 19 else
"1111111111111" when X = 56 AND Y = 19 else
"1111111111111" when X = 57 AND Y = 19 else
"1111111111111" when X = 58 AND Y = 19 else
"1111111111111" when X = 59 AND Y = 19 else
"1111111111111" when X = 60 AND Y = 19 else
"1111111111111" when X = 61 AND Y = 19 else
"1111111111111" when X = 62 AND Y = 19 else
"1101111011111" when X = 63 AND Y = 19 else
"1101110111111" when X = 64 AND Y = 19 else
"1100110011101" when X = 65 AND Y = 19 else
"1001101010111" when X = 66 AND Y = 19 else
"1001100110101" when X = 67 AND Y = 19 else
"0100010001001" when X = 68 AND Y = 19 else
"0000000000000" when X = 69 AND Y = 19 else
"0000000000000" when X = 70 AND Y = 19 else
"0000000000000" when X = 71 AND Y = 19 else
"0000000000000" when X = 72 AND Y = 19 else
"0000000000000" when X = 73 AND Y = 19 else
"0000000000000" when X = 74 AND Y = 19 else
"1000100111011" when X = 0 AND Y = 20 else
"1000100111011" when X = 1 AND Y = 20 else
"1000100111011" when X = 2 AND Y = 20 else
"1000100111011" when X = 3 AND Y = 20 else
"1000100111011" when X = 4 AND Y = 20 else
"1010101111101" when X = 5 AND Y = 20 else
"1101110111111" when X = 6 AND Y = 20 else
"1101110111111" when X = 7 AND Y = 20 else
"1101110111111" when X = 8 AND Y = 20 else
"1101110111111" when X = 9 AND Y = 20 else
"1101110111111" when X = 10 AND Y = 20 else
"1101110111111" when X = 11 AND Y = 20 else
"1101110111111" when X = 12 AND Y = 20 else
"1101110111111" when X = 13 AND Y = 20 else
"1101110111111" when X = 14 AND Y = 20 else
"1101110111111" when X = 15 AND Y = 20 else
"1110111011111" when X = 16 AND Y = 20 else
"1110111011111" when X = 17 AND Y = 20 else
"1110111011111" when X = 18 AND Y = 20 else
"1110111011111" when X = 19 AND Y = 20 else
"1110111011111" when X = 20 AND Y = 20 else
"1110111011111" when X = 21 AND Y = 20 else
"1110111011111" when X = 22 AND Y = 20 else
"1111111111111" when X = 23 AND Y = 20 else
"1111111111111" when X = 24 AND Y = 20 else
"1111111111111" when X = 25 AND Y = 20 else
"1111111111111" when X = 26 AND Y = 20 else
"1111111111111" when X = 27 AND Y = 20 else
"1111111111111" when X = 28 AND Y = 20 else
"1111111111111" when X = 29 AND Y = 20 else
"1111111111111" when X = 30 AND Y = 20 else
"1111111111111" when X = 31 AND Y = 20 else
"1111111111111" when X = 32 AND Y = 20 else
"1111111111111" when X = 33 AND Y = 20 else
"1111111111111" when X = 34 AND Y = 20 else
"1111111111111" when X = 35 AND Y = 20 else
"1111111111111" when X = 36 AND Y = 20 else
"1111111111111" when X = 37 AND Y = 20 else
"1111111111111" when X = 38 AND Y = 20 else
"1111111111111" when X = 39 AND Y = 20 else
"1111111111111" when X = 40 AND Y = 20 else
"1111111111111" when X = 41 AND Y = 20 else
"1111111111111" when X = 42 AND Y = 20 else
"1111111111111" when X = 43 AND Y = 20 else
"1111111111111" when X = 44 AND Y = 20 else
"1111111111111" when X = 45 AND Y = 20 else
"1111111111111" when X = 46 AND Y = 20 else
"1111111111111" when X = 47 AND Y = 20 else
"1111111111111" when X = 48 AND Y = 20 else
"1111111111111" when X = 49 AND Y = 20 else
"1111111111111" when X = 50 AND Y = 20 else
"1111111111111" when X = 51 AND Y = 20 else
"1111111111111" when X = 52 AND Y = 20 else
"1111111111111" when X = 53 AND Y = 20 else
"1111111111111" when X = 54 AND Y = 20 else
"1111111111111" when X = 55 AND Y = 20 else
"1111111111111" when X = 56 AND Y = 20 else
"1111111111111" when X = 57 AND Y = 20 else
"1111111111111" when X = 58 AND Y = 20 else
"1111111111111" when X = 59 AND Y = 20 else
"1111111111111" when X = 60 AND Y = 20 else
"1111111111111" when X = 61 AND Y = 20 else
"1111111111111" when X = 62 AND Y = 20 else
"1110111011111" when X = 63 AND Y = 20 else
"1101110111111" when X = 64 AND Y = 20 else
"1101110111111" when X = 65 AND Y = 20 else
"1101110111111" when X = 66 AND Y = 20 else
"1100110111101" when X = 67 AND Y = 20 else
"0101010101101" when X = 68 AND Y = 20 else
"0000000000000" when X = 69 AND Y = 20 else
"0000000000000" when X = 70 AND Y = 20 else
"0000000000000" when X = 71 AND Y = 20 else
"0000000000000" when X = 72 AND Y = 20 else
"0000000000000" when X = 73 AND Y = 20 else
"0000000000000" when X = 74 AND Y = 20 else
"1000100111011" when X = 0 AND Y = 21 else
"1000100111011" when X = 1 AND Y = 21 else
"1000100111011" when X = 2 AND Y = 21 else
"1000100111011" when X = 3 AND Y = 21 else
"1011101111101" when X = 4 AND Y = 21 else
"1101110111111" when X = 5 AND Y = 21 else
"1101110111111" when X = 6 AND Y = 21 else
"1101110111111" when X = 7 AND Y = 21 else
"1101110111111" when X = 8 AND Y = 21 else
"1101110111111" when X = 9 AND Y = 21 else
"1101110111111" when X = 10 AND Y = 21 else
"1101110111111" when X = 11 AND Y = 21 else
"1101110111111" when X = 12 AND Y = 21 else
"1101110111111" when X = 13 AND Y = 21 else
"1101110111111" when X = 14 AND Y = 21 else
"1101110111111" when X = 15 AND Y = 21 else
"1111111111111" when X = 16 AND Y = 21 else
"1111111111111" when X = 17 AND Y = 21 else
"1111111111111" when X = 18 AND Y = 21 else
"1111111111111" when X = 19 AND Y = 21 else
"1111111111111" when X = 20 AND Y = 21 else
"1111111111111" when X = 21 AND Y = 21 else
"1111111111111" when X = 22 AND Y = 21 else
"1111111111111" when X = 23 AND Y = 21 else
"1111111111111" when X = 24 AND Y = 21 else
"1111111111111" when X = 25 AND Y = 21 else
"1111111111111" when X = 26 AND Y = 21 else
"1111111111111" when X = 27 AND Y = 21 else
"1111111111111" when X = 28 AND Y = 21 else
"1111111111111" when X = 29 AND Y = 21 else
"1111111111111" when X = 30 AND Y = 21 else
"1111111111111" when X = 31 AND Y = 21 else
"1111111111111" when X = 32 AND Y = 21 else
"1111111111111" when X = 33 AND Y = 21 else
"1111111111111" when X = 34 AND Y = 21 else
"1111111111111" when X = 35 AND Y = 21 else
"1111111111111" when X = 36 AND Y = 21 else
"1111111111111" when X = 37 AND Y = 21 else
"1111111111111" when X = 38 AND Y = 21 else
"1111111111111" when X = 39 AND Y = 21 else
"1111111111111" when X = 40 AND Y = 21 else
"1111111111111" when X = 41 AND Y = 21 else
"1111111111111" when X = 42 AND Y = 21 else
"1111111111111" when X = 43 AND Y = 21 else
"1111111111111" when X = 44 AND Y = 21 else
"1111111111111" when X = 45 AND Y = 21 else
"1111111111111" when X = 46 AND Y = 21 else
"1111111111111" when X = 47 AND Y = 21 else
"1111111111111" when X = 48 AND Y = 21 else
"1111111111111" when X = 49 AND Y = 21 else
"1110111111111" when X = 50 AND Y = 21 else
"1110111011111" when X = 51 AND Y = 21 else
"1110111011111" when X = 52 AND Y = 21 else
"1111111111111" when X = 53 AND Y = 21 else
"1111111111111" when X = 54 AND Y = 21 else
"1111111111111" when X = 55 AND Y = 21 else
"1111111111111" when X = 56 AND Y = 21 else
"1111111111111" when X = 57 AND Y = 21 else
"1111111111111" when X = 58 AND Y = 21 else
"1111111111111" when X = 59 AND Y = 21 else
"1111111111111" when X = 60 AND Y = 21 else
"1111111111111" when X = 61 AND Y = 21 else
"1111111111111" when X = 62 AND Y = 21 else
"1110111011111" when X = 63 AND Y = 21 else
"1101110111111" when X = 64 AND Y = 21 else
"1101110111111" when X = 65 AND Y = 21 else
"1101111011111" when X = 66 AND Y = 21 else
"1101110111101" when X = 67 AND Y = 21 else
"1001100110011" when X = 68 AND Y = 21 else
"1000100010001" when X = 69 AND Y = 21 else
"0111011110001" when X = 70 AND Y = 21 else
"0110011101111" when X = 71 AND Y = 21 else
"0110011101111" when X = 72 AND Y = 21 else
"0110011101111" when X = 73 AND Y = 21 else
"0110011101111" when X = 74 AND Y = 21 else
"0111100011001" when X = 0 AND Y = 22 else
"1000100111011" when X = 1 AND Y = 22 else
"1000100111011" when X = 2 AND Y = 22 else
"1010101111101" when X = 3 AND Y = 22 else
"1100110111101" when X = 4 AND Y = 22 else
"1101110111111" when X = 5 AND Y = 22 else
"1101110111111" when X = 6 AND Y = 22 else
"1101110111111" when X = 7 AND Y = 22 else
"1101110111111" when X = 8 AND Y = 22 else
"1101110111111" when X = 9 AND Y = 22 else
"1101110111111" when X = 10 AND Y = 22 else
"1101110111111" when X = 11 AND Y = 22 else
"1101110111111" when X = 12 AND Y = 22 else
"1101110111111" when X = 13 AND Y = 22 else
"1101110111111" when X = 14 AND Y = 22 else
"1101110111111" when X = 15 AND Y = 22 else
"1111111111111" when X = 16 AND Y = 22 else
"1111111111111" when X = 17 AND Y = 22 else
"1111111111111" when X = 18 AND Y = 22 else
"1111111111111" when X = 19 AND Y = 22 else
"1111111111111" when X = 20 AND Y = 22 else
"1111111111111" when X = 21 AND Y = 22 else
"1111111111111" when X = 22 AND Y = 22 else
"1111111111111" when X = 23 AND Y = 22 else
"1111111111111" when X = 24 AND Y = 22 else
"1111111111111" when X = 25 AND Y = 22 else
"1111111111111" when X = 26 AND Y = 22 else
"1111111111111" when X = 27 AND Y = 22 else
"1111111111111" when X = 28 AND Y = 22 else
"1111111111111" when X = 29 AND Y = 22 else
"1111111111111" when X = 30 AND Y = 22 else
"1111111111111" when X = 31 AND Y = 22 else
"1111111111111" when X = 32 AND Y = 22 else
"1111111111111" when X = 33 AND Y = 22 else
"1111111111111" when X = 34 AND Y = 22 else
"1111111111111" when X = 35 AND Y = 22 else
"1111111111111" when X = 36 AND Y = 22 else
"1111111111111" when X = 37 AND Y = 22 else
"1111111111111" when X = 38 AND Y = 22 else
"1111111111111" when X = 39 AND Y = 22 else
"1111111111111" when X = 40 AND Y = 22 else
"1111111111111" when X = 41 AND Y = 22 else
"1111111111111" when X = 42 AND Y = 22 else
"1111111111111" when X = 43 AND Y = 22 else
"1111111111111" when X = 44 AND Y = 22 else
"1111111111111" when X = 45 AND Y = 22 else
"1111111111111" when X = 46 AND Y = 22 else
"1110111011111" when X = 47 AND Y = 22 else
"1101110111111" when X = 48 AND Y = 22 else
"1101110111111" when X = 49 AND Y = 22 else
"1110111011111" when X = 50 AND Y = 22 else
"1111111111111" when X = 51 AND Y = 22 else
"1111111111111" when X = 52 AND Y = 22 else
"1111111111111" when X = 53 AND Y = 22 else
"1111111111111" when X = 54 AND Y = 22 else
"1111111111111" when X = 55 AND Y = 22 else
"1111111111111" when X = 56 AND Y = 22 else
"1111111111111" when X = 57 AND Y = 22 else
"1111111111111" when X = 58 AND Y = 22 else
"1111111111111" when X = 59 AND Y = 22 else
"1111111111111" when X = 60 AND Y = 22 else
"1111111111111" when X = 61 AND Y = 22 else
"1111111111111" when X = 62 AND Y = 22 else
"1110111011111" when X = 63 AND Y = 22 else
"1101110111111" when X = 64 AND Y = 22 else
"1110111011111" when X = 65 AND Y = 22 else
"1111111111111" when X = 66 AND Y = 22 else
"1111111111111" when X = 67 AND Y = 22 else
"1111111111111" when X = 68 AND Y = 22 else
"1111111111111" when X = 69 AND Y = 22 else
"1110111011111" when X = 70 AND Y = 22 else
"1101110111101" when X = 71 AND Y = 22 else
"1101110111101" when X = 72 AND Y = 22 else
"1101110111101" when X = 73 AND Y = 22 else
"1101110111101" when X = 74 AND Y = 22 else
"0011001101011" when X = 0 AND Y = 23 else
"0111100011001" when X = 1 AND Y = 23 else
"1000100111011" when X = 2 AND Y = 23 else
"1000100111011" when X = 3 AND Y = 23 else
"1010101111101" when X = 4 AND Y = 23 else
"1101110111111" when X = 5 AND Y = 23 else
"1101110111111" when X = 6 AND Y = 23 else
"1101110111111" when X = 7 AND Y = 23 else
"1101110111111" when X = 8 AND Y = 23 else
"1101110111111" when X = 9 AND Y = 23 else
"1101110111111" when X = 10 AND Y = 23 else
"1101110111111" when X = 11 AND Y = 23 else
"1101110111111" when X = 12 AND Y = 23 else
"1101110111111" when X = 13 AND Y = 23 else
"1101110111111" when X = 14 AND Y = 23 else
"1101110111111" when X = 15 AND Y = 23 else
"1111111111111" when X = 16 AND Y = 23 else
"1111111111111" when X = 17 AND Y = 23 else
"1111111111111" when X = 18 AND Y = 23 else
"1111111111111" when X = 19 AND Y = 23 else
"1111111111111" when X = 20 AND Y = 23 else
"1111111111111" when X = 21 AND Y = 23 else
"1111111111111" when X = 22 AND Y = 23 else
"1111111111111" when X = 23 AND Y = 23 else
"1111111111111" when X = 24 AND Y = 23 else
"1111111111111" when X = 25 AND Y = 23 else
"1111111111111" when X = 26 AND Y = 23 else
"1111111111111" when X = 27 AND Y = 23 else
"1111111111111" when X = 28 AND Y = 23 else
"1111111111111" when X = 29 AND Y = 23 else
"1111111111111" when X = 30 AND Y = 23 else
"1111111111111" when X = 31 AND Y = 23 else
"1111111111111" when X = 32 AND Y = 23 else
"1111111111111" when X = 33 AND Y = 23 else
"1111111111111" when X = 34 AND Y = 23 else
"1111111111111" when X = 35 AND Y = 23 else
"1111111111111" when X = 36 AND Y = 23 else
"1101111011111" when X = 37 AND Y = 23 else
"1101110111111" when X = 38 AND Y = 23 else
"1101110111111" when X = 39 AND Y = 23 else
"1101110111111" when X = 40 AND Y = 23 else
"1101110111111" when X = 41 AND Y = 23 else
"1101110111111" when X = 42 AND Y = 23 else
"1101110111111" when X = 43 AND Y = 23 else
"1101110111111" when X = 44 AND Y = 23 else
"1101110111111" when X = 45 AND Y = 23 else
"1101110111111" when X = 46 AND Y = 23 else
"1101110111111" when X = 47 AND Y = 23 else
"1101110111111" when X = 48 AND Y = 23 else
"1110111011111" when X = 49 AND Y = 23 else
"1111111111111" when X = 50 AND Y = 23 else
"1111111111111" when X = 51 AND Y = 23 else
"1111111111111" when X = 52 AND Y = 23 else
"1111111111111" when X = 53 AND Y = 23 else
"1111111111111" when X = 54 AND Y = 23 else
"1110111011111" when X = 55 AND Y = 23 else
"1101110111101" when X = 56 AND Y = 23 else
"1110111011111" when X = 57 AND Y = 23 else
"1111111111111" when X = 58 AND Y = 23 else
"1111111111111" when X = 59 AND Y = 23 else
"1111111111111" when X = 60 AND Y = 23 else
"1111111111111" when X = 61 AND Y = 23 else
"1111111111111" when X = 62 AND Y = 23 else
"1110111011111" when X = 63 AND Y = 23 else
"1110111011111" when X = 64 AND Y = 23 else
"1111111111111" when X = 65 AND Y = 23 else
"1111111111111" when X = 66 AND Y = 23 else
"1111111111111" when X = 67 AND Y = 23 else
"1111111111111" when X = 68 AND Y = 23 else
"1111111111111" when X = 69 AND Y = 23 else
"1110111011111" when X = 70 AND Y = 23 else
"1101110111111" when X = 71 AND Y = 23 else
"1101110111111" when X = 72 AND Y = 23 else
"1101110111111" when X = 73 AND Y = 23 else
"1101110111111" when X = 74 AND Y = 23 else
"0001000100111" when X = 0 AND Y = 24 else
"0111100011001" when X = 1 AND Y = 24 else
"1000100111011" when X = 2 AND Y = 24 else
"1000100111011" when X = 3 AND Y = 24 else
"1000100111011" when X = 4 AND Y = 24 else
"1010101111101" when X = 5 AND Y = 24 else
"1101110111111" when X = 6 AND Y = 24 else
"1101110111111" when X = 7 AND Y = 24 else
"1101110111111" when X = 8 AND Y = 24 else
"1101110111111" when X = 9 AND Y = 24 else
"1101110111111" when X = 10 AND Y = 24 else
"1101110111111" when X = 11 AND Y = 24 else
"1101110111111" when X = 12 AND Y = 24 else
"1101110111111" when X = 13 AND Y = 24 else
"1101110111111" when X = 14 AND Y = 24 else
"1101110111111" when X = 15 AND Y = 24 else
"1111111111111" when X = 16 AND Y = 24 else
"1111111111111" when X = 17 AND Y = 24 else
"1111111111111" when X = 18 AND Y = 24 else
"1111111111111" when X = 19 AND Y = 24 else
"1111111111111" when X = 20 AND Y = 24 else
"1111111111111" when X = 21 AND Y = 24 else
"1111111111111" when X = 22 AND Y = 24 else
"1111111111111" when X = 23 AND Y = 24 else
"1111111111111" when X = 24 AND Y = 24 else
"1111111111111" when X = 25 AND Y = 24 else
"1111111111111" when X = 26 AND Y = 24 else
"1111111111111" when X = 27 AND Y = 24 else
"1111111111111" when X = 28 AND Y = 24 else
"1111111111111" when X = 29 AND Y = 24 else
"1111111111111" when X = 30 AND Y = 24 else
"1111111111111" when X = 31 AND Y = 24 else
"1111111111111" when X = 32 AND Y = 24 else
"1111111111111" when X = 33 AND Y = 24 else
"1111111111111" when X = 34 AND Y = 24 else
"1111111111111" when X = 35 AND Y = 24 else
"1111111111111" when X = 36 AND Y = 24 else
"1101110111111" when X = 37 AND Y = 24 else
"1101110111111" when X = 38 AND Y = 24 else
"1101110111111" when X = 39 AND Y = 24 else
"1101110111111" when X = 40 AND Y = 24 else
"1101110111111" when X = 41 AND Y = 24 else
"1101110111111" when X = 42 AND Y = 24 else
"1101110111111" when X = 43 AND Y = 24 else
"1101110111111" when X = 44 AND Y = 24 else
"1101110111111" when X = 45 AND Y = 24 else
"1101110111111" when X = 46 AND Y = 24 else
"1110111011111" when X = 47 AND Y = 24 else
"1111111111111" when X = 48 AND Y = 24 else
"1110111011111" when X = 49 AND Y = 24 else
"1101111011111" when X = 50 AND Y = 24 else
"1101111011111" when X = 51 AND Y = 24 else
"1101111011111" when X = 52 AND Y = 24 else
"1101111011111" when X = 53 AND Y = 24 else
"1101111011111" when X = 54 AND Y = 24 else
"1101110111111" when X = 55 AND Y = 24 else
"1010101011001" when X = 56 AND Y = 24 else
"1001100110101" when X = 57 AND Y = 24 else
"1101111011111" when X = 58 AND Y = 24 else
"1101111011111" when X = 59 AND Y = 24 else
"1101111011111" when X = 60 AND Y = 24 else
"1101111011111" when X = 61 AND Y = 24 else
"1101111011111" when X = 62 AND Y = 24 else
"1101110111111" when X = 63 AND Y = 24 else
"1110111011111" when X = 64 AND Y = 24 else
"1111111111111" when X = 65 AND Y = 24 else
"1111111111111" when X = 66 AND Y = 24 else
"1111111111111" when X = 67 AND Y = 24 else
"1111111111111" when X = 68 AND Y = 24 else
"1111111111111" when X = 69 AND Y = 24 else
"1110111011111" when X = 70 AND Y = 24 else
"1101110111111" when X = 71 AND Y = 24 else
"1101110111111" when X = 72 AND Y = 24 else
"1101110111111" when X = 73 AND Y = 24 else
"1101110111111" when X = 74 AND Y = 24 else
"0000000000011" when X = 0 AND Y = 25 else
"0100010001111" when X = 1 AND Y = 25 else
"0111100011001" when X = 2 AND Y = 25 else
"1000100111011" when X = 3 AND Y = 25 else
"1000100111011" when X = 4 AND Y = 25 else
"1001101011101" when X = 5 AND Y = 25 else
"1101110111111" when X = 6 AND Y = 25 else
"1101110111111" when X = 7 AND Y = 25 else
"1101110111111" when X = 8 AND Y = 25 else
"1101110111111" when X = 9 AND Y = 25 else
"1101110111111" when X = 10 AND Y = 25 else
"1101110111111" when X = 11 AND Y = 25 else
"1101110111111" when X = 12 AND Y = 25 else
"1101110111111" when X = 13 AND Y = 25 else
"1101110111111" when X = 14 AND Y = 25 else
"1101110111111" when X = 15 AND Y = 25 else
"1111111111111" when X = 16 AND Y = 25 else
"1111111111111" when X = 17 AND Y = 25 else
"1111111111111" when X = 18 AND Y = 25 else
"1111111111111" when X = 19 AND Y = 25 else
"1111111111111" when X = 20 AND Y = 25 else
"1111111111111" when X = 21 AND Y = 25 else
"1111111111111" when X = 22 AND Y = 25 else
"1111111111111" when X = 23 AND Y = 25 else
"1111111111111" when X = 24 AND Y = 25 else
"1111111111111" when X = 25 AND Y = 25 else
"1111111111111" when X = 26 AND Y = 25 else
"1111111111111" when X = 27 AND Y = 25 else
"1111111111111" when X = 28 AND Y = 25 else
"1111111111111" when X = 29 AND Y = 25 else
"1111111111111" when X = 30 AND Y = 25 else
"1111111111111" when X = 31 AND Y = 25 else
"1111111111111" when X = 32 AND Y = 25 else
"1111111111111" when X = 33 AND Y = 25 else
"1111111111111" when X = 34 AND Y = 25 else
"1111111111111" when X = 35 AND Y = 25 else
"1111111111111" when X = 36 AND Y = 25 else
"1111111111111" when X = 37 AND Y = 25 else
"1111111111111" when X = 38 AND Y = 25 else
"1111111111111" when X = 39 AND Y = 25 else
"1111111111111" when X = 40 AND Y = 25 else
"1111111111111" when X = 41 AND Y = 25 else
"1111111111111" when X = 42 AND Y = 25 else
"1111111111111" when X = 43 AND Y = 25 else
"1111111111111" when X = 44 AND Y = 25 else
"1111111111111" when X = 45 AND Y = 25 else
"1111111111111" when X = 46 AND Y = 25 else
"1111111111111" when X = 47 AND Y = 25 else
"1111111111111" when X = 48 AND Y = 25 else
"1101111011111" when X = 49 AND Y = 25 else
"1100110011011" when X = 50 AND Y = 25 else
"0111100010001" when X = 51 AND Y = 25 else
"0111011110001" when X = 52 AND Y = 25 else
"0111011110001" when X = 53 AND Y = 25 else
"0111011110001" when X = 54 AND Y = 25 else
"0111011110001" when X = 55 AND Y = 25 else
"0101010101101" when X = 56 AND Y = 25 else
"0111100010011" when X = 57 AND Y = 25 else
"1101110111111" when X = 58 AND Y = 25 else
"1101110111111" when X = 59 AND Y = 25 else
"1101110111111" when X = 60 AND Y = 25 else
"1101110111111" when X = 61 AND Y = 25 else
"1101110111111" when X = 62 AND Y = 25 else
"1101110111111" when X = 63 AND Y = 25 else
"1110111011111" when X = 64 AND Y = 25 else
"1111111111111" when X = 65 AND Y = 25 else
"1111111111111" when X = 66 AND Y = 25 else
"1111111111111" when X = 67 AND Y = 25 else
"1111111111111" when X = 68 AND Y = 25 else
"1111111111111" when X = 69 AND Y = 25 else
"1110111011111" when X = 70 AND Y = 25 else
"1101110111111" when X = 71 AND Y = 25 else
"1101110111111" when X = 72 AND Y = 25 else
"1101110111111" when X = 73 AND Y = 25 else
"1101110111111" when X = 74 AND Y = 25 else
"0000000000000" when X = 0 AND Y = 26 else
"0000000000000" when X = 1 AND Y = 26 else
"0110011110111" when X = 2 AND Y = 26 else
"1000100111011" when X = 3 AND Y = 26 else
"1000100111011" when X = 4 AND Y = 26 else
"1000100111011" when X = 5 AND Y = 26 else
"1010101111101" when X = 6 AND Y = 26 else
"1101110111111" when X = 7 AND Y = 26 else
"1101110111111" when X = 8 AND Y = 26 else
"1101110111111" when X = 9 AND Y = 26 else
"1101110111111" when X = 10 AND Y = 26 else
"1101110111111" when X = 11 AND Y = 26 else
"1101110111111" when X = 12 AND Y = 26 else
"1101110111111" when X = 13 AND Y = 26 else
"1101110111111" when X = 14 AND Y = 26 else
"1101110111111" when X = 15 AND Y = 26 else
"1110111011111" when X = 16 AND Y = 26 else
"1110111011111" when X = 17 AND Y = 26 else
"1110111011111" when X = 18 AND Y = 26 else
"1110111011111" when X = 19 AND Y = 26 else
"1110111011111" when X = 20 AND Y = 26 else
"1110111011111" when X = 21 AND Y = 26 else
"1110111011111" when X = 22 AND Y = 26 else
"1110111011111" when X = 23 AND Y = 26 else
"1110111011111" when X = 24 AND Y = 26 else
"1110111011111" when X = 25 AND Y = 26 else
"1110111011111" when X = 26 AND Y = 26 else
"1110111011111" when X = 27 AND Y = 26 else
"1110111011111" when X = 28 AND Y = 26 else
"1110111011111" when X = 29 AND Y = 26 else
"1110111011111" when X = 30 AND Y = 26 else
"1110111011111" when X = 31 AND Y = 26 else
"1110111011111" when X = 32 AND Y = 26 else
"1111111111111" when X = 33 AND Y = 26 else
"1111111111111" when X = 34 AND Y = 26 else
"1111111111111" when X = 35 AND Y = 26 else
"1111111111111" when X = 36 AND Y = 26 else
"1111111111111" when X = 37 AND Y = 26 else
"1111111111111" when X = 38 AND Y = 26 else
"1111111111111" when X = 39 AND Y = 26 else
"1111111111111" when X = 40 AND Y = 26 else
"1111111111111" when X = 41 AND Y = 26 else
"1111111111111" when X = 42 AND Y = 26 else
"1111111111111" when X = 43 AND Y = 26 else
"1111111111111" when X = 44 AND Y = 26 else
"1111111111111" when X = 45 AND Y = 26 else
"1111111111111" when X = 46 AND Y = 26 else
"1111111111111" when X = 47 AND Y = 26 else
"1101111011111" when X = 48 AND Y = 26 else
"1101110111111" when X = 49 AND Y = 26 else
"1011101111011" when X = 50 AND Y = 26 else
"0001000100011" when X = 51 AND Y = 26 else
"0000000000000" when X = 52 AND Y = 26 else
"0000000000000" when X = 53 AND Y = 26 else
"0000000000000" when X = 54 AND Y = 26 else
"0000000000000" when X = 55 AND Y = 26 else
"0000000000000" when X = 56 AND Y = 26 else
"1000100010011" when X = 57 AND Y = 26 else
"1101110111111" when X = 58 AND Y = 26 else
"1101110111111" when X = 59 AND Y = 26 else
"1101110111111" when X = 60 AND Y = 26 else
"1101110111111" when X = 61 AND Y = 26 else
"1101110111111" when X = 62 AND Y = 26 else
"1101110111111" when X = 63 AND Y = 26 else
"1110111011111" when X = 64 AND Y = 26 else
"1111111111111" when X = 65 AND Y = 26 else
"1111111111111" when X = 66 AND Y = 26 else
"1111111111111" when X = 67 AND Y = 26 else
"1111111111111" when X = 68 AND Y = 26 else
"1110111111111" when X = 69 AND Y = 26 else
"1101111011111" when X = 70 AND Y = 26 else
"1101110111111" when X = 71 AND Y = 26 else
"1101110111111" when X = 72 AND Y = 26 else
"1101110111111" when X = 73 AND Y = 26 else
"1101110111111" when X = 74 AND Y = 26 else
"0000000000000" when X = 0 AND Y = 27 else
"0000000000001" when X = 1 AND Y = 27 else
"0101010110001" when X = 2 AND Y = 27 else
"0110011010101" when X = 3 AND Y = 27 else
"0111100010111" when X = 4 AND Y = 27 else
"1000100111011" when X = 5 AND Y = 27 else
"1000100111011" when X = 6 AND Y = 27 else
"1010101111101" when X = 7 AND Y = 27 else
"1011101111101" when X = 8 AND Y = 27 else
"1100110111101" when X = 9 AND Y = 27 else
"1101110111111" when X = 10 AND Y = 27 else
"1101110111111" when X = 11 AND Y = 27 else
"1101110111111" when X = 12 AND Y = 27 else
"1101110111111" when X = 13 AND Y = 27 else
"1101110111111" when X = 14 AND Y = 27 else
"1101110111111" when X = 15 AND Y = 27 else
"1101110111111" when X = 16 AND Y = 27 else
"1101110111111" when X = 17 AND Y = 27 else
"1101110111111" when X = 18 AND Y = 27 else
"1101110111111" when X = 19 AND Y = 27 else
"1101110111111" when X = 20 AND Y = 27 else
"1101110111111" when X = 21 AND Y = 27 else
"1101110111111" when X = 22 AND Y = 27 else
"1101110111111" when X = 23 AND Y = 27 else
"1101110111111" when X = 24 AND Y = 27 else
"1101110111111" when X = 25 AND Y = 27 else
"1101110111111" when X = 26 AND Y = 27 else
"1101110111111" when X = 27 AND Y = 27 else
"1101110111111" when X = 28 AND Y = 27 else
"1101110111111" when X = 29 AND Y = 27 else
"1101110111111" when X = 30 AND Y = 27 else
"1101110111111" when X = 31 AND Y = 27 else
"1101110111111" when X = 32 AND Y = 27 else
"1110111011111" when X = 33 AND Y = 27 else
"1110111011111" when X = 34 AND Y = 27 else
"1110111011111" when X = 35 AND Y = 27 else
"1110111011111" when X = 36 AND Y = 27 else
"1110111111111" when X = 37 AND Y = 27 else
"1111111111111" when X = 38 AND Y = 27 else
"1111111111111" when X = 39 AND Y = 27 else
"1111111111111" when X = 40 AND Y = 27 else
"1111111111111" when X = 41 AND Y = 27 else
"1111111111111" when X = 42 AND Y = 27 else
"1111111111111" when X = 43 AND Y = 27 else
"1110111111111" when X = 44 AND Y = 27 else
"1110111011111" when X = 45 AND Y = 27 else
"1110111011111" when X = 46 AND Y = 27 else
"1101111011111" when X = 47 AND Y = 27 else
"1101110111111" when X = 48 AND Y = 27 else
"1101110111111" when X = 49 AND Y = 27 else
"1011110011011" when X = 50 AND Y = 27 else
"0010001000101" when X = 51 AND Y = 27 else
"0000000000000" when X = 52 AND Y = 27 else
"0000000000000" when X = 53 AND Y = 27 else
"0000000000000" when X = 54 AND Y = 27 else
"0000000000000" when X = 55 AND Y = 27 else
"0000000000000" when X = 56 AND Y = 27 else
"0110011001111" when X = 57 AND Y = 27 else
"1011101111001" when X = 58 AND Y = 27 else
"1101110111101" when X = 59 AND Y = 27 else
"1101110111111" when X = 60 AND Y = 27 else
"1101110111111" when X = 61 AND Y = 27 else
"1101110111111" when X = 62 AND Y = 27 else
"1101110111111" when X = 63 AND Y = 27 else
"1101111011111" when X = 64 AND Y = 27 else
"1110111011111" when X = 65 AND Y = 27 else
"1110111011111" when X = 66 AND Y = 27 else
"1110111011111" when X = 67 AND Y = 27 else
"1110111011111" when X = 68 AND Y = 27 else
"1101111011111" when X = 69 AND Y = 27 else
"1101110111111" when X = 70 AND Y = 27 else
"1101110111111" when X = 71 AND Y = 27 else
"1101110111111" when X = 72 AND Y = 27 else
"1101110111111" when X = 73 AND Y = 27 else
"1101110111111" when X = 74 AND Y = 27 else
"0000000000000" when X = 0 AND Y = 28 else
"0000000000000" when X = 1 AND Y = 28 else
"0000000000000" when X = 2 AND Y = 28 else
"0000000000000" when X = 3 AND Y = 28 else
"0100010001111" when X = 4 AND Y = 28 else
"0110011110111" when X = 5 AND Y = 28 else
"0111011110111" when X = 6 AND Y = 28 else
"1000100111011" when X = 7 AND Y = 28 else
"1000100111011" when X = 8 AND Y = 28 else
"1010101111101" when X = 9 AND Y = 28 else
"1011110011101" when X = 10 AND Y = 28 else
"1011110011101" when X = 11 AND Y = 28 else
"1011110011101" when X = 12 AND Y = 28 else
"1011110011101" when X = 13 AND Y = 28 else
"1011110011101" when X = 14 AND Y = 28 else
"1011110011101" when X = 15 AND Y = 28 else
"1011110011101" when X = 16 AND Y = 28 else
"1011110011101" when X = 17 AND Y = 28 else
"1011110011101" when X = 18 AND Y = 28 else
"1011110011101" when X = 19 AND Y = 28 else
"1011110011101" when X = 20 AND Y = 28 else
"1011110011101" when X = 21 AND Y = 28 else
"1011110011101" when X = 22 AND Y = 28 else
"1011101111011" when X = 23 AND Y = 28 else
"1011101111001" when X = 24 AND Y = 28 else
"1011101111001" when X = 25 AND Y = 28 else
"1011101111001" when X = 26 AND Y = 28 else
"1011101111001" when X = 27 AND Y = 28 else
"1011110011011" when X = 28 AND Y = 28 else
"1101110111111" when X = 29 AND Y = 28 else
"1101110111111" when X = 30 AND Y = 28 else
"1101110111111" when X = 31 AND Y = 28 else
"1101110111111" when X = 32 AND Y = 28 else
"1101110111111" when X = 33 AND Y = 28 else
"1101110111111" when X = 34 AND Y = 28 else
"1101110111111" when X = 35 AND Y = 28 else
"1101110111111" when X = 36 AND Y = 28 else
"1101110111111" when X = 37 AND Y = 28 else
"1110111011111" when X = 38 AND Y = 28 else
"1111111111111" when X = 39 AND Y = 28 else
"1111111111111" when X = 40 AND Y = 28 else
"1111111111111" when X = 41 AND Y = 28 else
"1111111111111" when X = 42 AND Y = 28 else
"1110111011111" when X = 43 AND Y = 28 else
"1101110111111" when X = 44 AND Y = 28 else
"1101110111111" when X = 45 AND Y = 28 else
"1101110111111" when X = 46 AND Y = 28 else
"1101110111111" when X = 47 AND Y = 28 else
"1101110111111" when X = 48 AND Y = 28 else
"1100110011101" when X = 49 AND Y = 28 else
"1001101010111" when X = 50 AND Y = 28 else
"0001000100011" when X = 51 AND Y = 28 else
"0000000000000" when X = 52 AND Y = 28 else
"0000000000000" when X = 53 AND Y = 28 else
"0000000000000" when X = 54 AND Y = 28 else
"0000000000000" when X = 55 AND Y = 28 else
"0000000000000" when X = 56 AND Y = 28 else
"0000000000000" when X = 57 AND Y = 28 else
"0110011001111" when X = 58 AND Y = 28 else
"1101110111101" when X = 59 AND Y = 28 else
"1101110111111" when X = 60 AND Y = 28 else
"1101110111111" when X = 61 AND Y = 28 else
"1101110111111" when X = 62 AND Y = 28 else
"1101110111111" when X = 63 AND Y = 28 else
"1101110111111" when X = 64 AND Y = 28 else
"1100110111101" when X = 65 AND Y = 28 else
"1011101111001" when X = 66 AND Y = 28 else
"1011101111001" when X = 67 AND Y = 28 else
"1011101111001" when X = 68 AND Y = 28 else
"1011101111001" when X = 69 AND Y = 28 else
"1011101111001" when X = 70 AND Y = 28 else
"1011101111001" when X = 71 AND Y = 28 else
"1011101111001" when X = 72 AND Y = 28 else
"1011101111001" when X = 73 AND Y = 28 else
"1011101111001" when X = 74 AND Y = 28 else
"0000000000000" when X = 0 AND Y = 29 else
"0000000000000" when X = 1 AND Y = 29 else
"0000000000000" when X = 2 AND Y = 29 else
"0000000000000" when X = 3 AND Y = 29 else
"0000000000001" when X = 4 AND Y = 29 else
"0000000000011" when X = 5 AND Y = 29 else
"0011001101011" when X = 6 AND Y = 29 else
"0111011110111" when X = 7 AND Y = 29 else
"0111100011001" when X = 8 AND Y = 29 else
"1000100111011" when X = 9 AND Y = 29 else
"1000100111011" when X = 10 AND Y = 29 else
"1000100111011" when X = 11 AND Y = 29 else
"1000100111011" when X = 12 AND Y = 29 else
"1000100111011" when X = 13 AND Y = 29 else
"1000100111011" when X = 14 AND Y = 29 else
"1000100111011" when X = 15 AND Y = 29 else
"1000100111011" when X = 16 AND Y = 29 else
"1000100111011" when X = 17 AND Y = 29 else
"1000100111011" when X = 18 AND Y = 29 else
"0111100011011" when X = 19 AND Y = 29 else
"0111100011001" when X = 20 AND Y = 29 else
"0111100011001" when X = 21 AND Y = 29 else
"0111011110111" when X = 22 AND Y = 29 else
"0011001101011" when X = 23 AND Y = 29 else
"0001000100011" when X = 24 AND Y = 29 else
"0001000100011" when X = 25 AND Y = 29 else
"0001000100011" when X = 26 AND Y = 29 else
"0001000100011" when X = 27 AND Y = 29 else
"0110011001101" when X = 28 AND Y = 29 else
"1011110011011" when X = 29 AND Y = 29 else
"1100110011011" when X = 30 AND Y = 29 else
"1101110111101" when X = 31 AND Y = 29 else
"1101110111111" when X = 32 AND Y = 29 else
"1101110111111" when X = 33 AND Y = 29 else
"1101110111111" when X = 34 AND Y = 29 else
"1101110111111" when X = 35 AND Y = 29 else
"1101110111111" when X = 36 AND Y = 29 else
"1101110111111" when X = 37 AND Y = 29 else
"1101110111111" when X = 38 AND Y = 29 else
"1101110111111" when X = 39 AND Y = 29 else
"1101110111111" when X = 40 AND Y = 29 else
"1101110111111" when X = 41 AND Y = 29 else
"1101110111111" when X = 42 AND Y = 29 else
"1101110111111" when X = 43 AND Y = 29 else
"1101110111101" when X = 44 AND Y = 29 else
"1100110011011" when X = 45 AND Y = 29 else
"1100110011011" when X = 46 AND Y = 29 else
"1100110011011" when X = 47 AND Y = 29 else
"1100110011011" when X = 48 AND Y = 29 else
"1001100110101" when X = 49 AND Y = 29 else
"0001000100011" when X = 50 AND Y = 29 else
"0000000000000" when X = 51 AND Y = 29 else
"0000000000000" when X = 52 AND Y = 29 else
"0000000000000" when X = 53 AND Y = 29 else
"0000000000000" when X = 54 AND Y = 29 else
"0000000000000" when X = 55 AND Y = 29 else
"0000000000000" when X = 56 AND Y = 29 else
"0000000000000" when X = 57 AND Y = 29 else
"0101011001101" when X = 58 AND Y = 29 else
"1011110011011" when X = 59 AND Y = 29 else
"1100110011011" when X = 60 AND Y = 29 else
"1100110011011" when X = 61 AND Y = 29 else
"1100110011011" when X = 62 AND Y = 29 else
"1100110011011" when X = 63 AND Y = 29 else
"1100110011011" when X = 64 AND Y = 29 else
"1010101010111" when X = 65 AND Y = 29 else
"0010001000101" when X = 66 AND Y = 29 else
"0001000100011" when X = 67 AND Y = 29 else
"0001000100011" when X = 68 AND Y = 29 else
"0001000100011" when X = 69 AND Y = 29 else
"0001000100011" when X = 70 AND Y = 29 else
"0001000100011" when X = 71 AND Y = 29 else
"0001000100011" when X = 72 AND Y = 29 else
"0001000100011" when X = 73 AND Y = 29 else
"0001000100011" when X = 74 AND Y = 29 else
"0000000000000" when X = 0 AND Y = 30 else
"0000000000000" when X = 1 AND Y = 30 else
"0000000000000" when X = 2 AND Y = 30 else
"0000000000000" when X = 3 AND Y = 30 else
"0000000000000" when X = 4 AND Y = 30 else
"0000000000000" when X = 5 AND Y = 30 else
"0000000000011" when X = 6 AND Y = 30 else
"0001001000111" when X = 7 AND Y = 30 else
"0010001001001" when X = 8 AND Y = 30 else
"0111100010111" when X = 9 AND Y = 30 else
"1000100111011" when X = 10 AND Y = 30 else
"1000100111011" when X = 11 AND Y = 30 else
"1000100111011" when X = 12 AND Y = 30 else
"1000100111011" when X = 13 AND Y = 30 else
"1000100111011" when X = 14 AND Y = 30 else
"1000100111011" when X = 15 AND Y = 30 else
"1000100111011" when X = 16 AND Y = 30 else
"1000100111011" when X = 17 AND Y = 30 else
"1000100111011" when X = 18 AND Y = 30 else
"0110011110111" when X = 19 AND Y = 30 else
"0001001000111" when X = 20 AND Y = 30 else
"0001001000111" when X = 21 AND Y = 30 else
"0001001000111" when X = 22 AND Y = 30 else
"0000000000011" when X = 23 AND Y = 30 else
"0000000000000" when X = 24 AND Y = 30 else
"0000000000000" when X = 25 AND Y = 30 else
"0000000000000" when X = 26 AND Y = 30 else
"0000000000000" when X = 27 AND Y = 30 else
"0001000100011" when X = 28 AND Y = 30 else
"0011001100111" when X = 29 AND Y = 30 else
"0100010001011" when X = 30 AND Y = 30 else
"1100110011011" when X = 31 AND Y = 30 else
"1101110111111" when X = 32 AND Y = 30 else
"1101110111111" when X = 33 AND Y = 30 else
"1101110111111" when X = 34 AND Y = 30 else
"1101110111111" when X = 35 AND Y = 30 else
"1101110111111" when X = 36 AND Y = 30 else
"1101110111111" when X = 37 AND Y = 30 else
"1101110111111" when X = 38 AND Y = 30 else
"1101110111111" when X = 39 AND Y = 30 else
"1101110111111" when X = 40 AND Y = 30 else
"1101110111111" when X = 41 AND Y = 30 else
"1101110111111" when X = 42 AND Y = 30 else
"1101110111111" when X = 43 AND Y = 30 else
"1100110111101" when X = 44 AND Y = 30 else
"0101011001101" when X = 45 AND Y = 30 else
"0011001101001" when X = 46 AND Y = 30 else
"0011001101001" when X = 47 AND Y = 30 else
"0011001101001" when X = 48 AND Y = 30 else
"0010001000111" when X = 49 AND Y = 30 else
"0000000000000" when X = 50 AND Y = 30 else
"0000000000000" when X = 51 AND Y = 30 else
"0000000000000" when X = 52 AND Y = 30 else
"0000000000000" when X = 53 AND Y = 30 else
"0000000000000" when X = 54 AND Y = 30 else
"0000000000000" when X = 55 AND Y = 30 else
"0000000000000" when X = 56 AND Y = 30 else
"0000000000000" when X = 57 AND Y = 30 else
"0001000100011" when X = 58 AND Y = 30 else
"0011001100111" when X = 59 AND Y = 30 else
"0011001101001" when X = 60 AND Y = 30 else
"0011001101001" when X = 61 AND Y = 30 else
"0011001101001" when X = 62 AND Y = 30 else
"0011001101001" when X = 63 AND Y = 30 else
"0011001101001" when X = 64 AND Y = 30 else
"0011001100111" when X = 65 AND Y = 30 else
"0000000000000" when X = 66 AND Y = 30 else
"0000000000000" when X = 67 AND Y = 30 else
"0000000000000" when X = 68 AND Y = 30 else
"0000000000000" when X = 69 AND Y = 30 else
"0000000000000" when X = 70 AND Y = 30 else
"0000000000000" when X = 71 AND Y = 30 else
"0000000000000" when X = 72 AND Y = 30 else
"0000000000000" when X = 73 AND Y = 30 else
"0000000000000" when X = 74 AND Y = 30 else
"0000000000000"; -- should never get here
end rtl;
