-- Tyler Hansen
-- CS232 Final Project
-- genSpriteROM.py
-- generates a ROM file in VHDL from a .ppm image

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity player_sprite_straight_updated is
port(
X	: in INTEGER RANGE 0 TO 1688;
Y	: in INTEGER RANGE 0 TO 1688;
data : out std_logic_vector (12 downto 0)
);

end entity;

architecture rtl of player_sprite_straight_updated is
begin
data <=
"1111111100000" when X = 0 AND Y = 0 else
"1111111100000" when X = 1 AND Y = 0 else
"1111111100000" when X = 2 AND Y = 0 else
"1111111100000" when X = 3 AND Y = 0 else
"1111111100000" when X = 4 AND Y = 0 else
"1111111100000" when X = 5 AND Y = 0 else
"1111111100000" when X = 6 AND Y = 0 else
"1111111100000" when X = 7 AND Y = 0 else
"1111111100000" when X = 8 AND Y = 0 else
"1111111100000" when X = 9 AND Y = 0 else
"1111111100000" when X = 10 AND Y = 0 else
"1111111100000" when X = 11 AND Y = 0 else
"1111111100000" when X = 12 AND Y = 0 else
"1111111100000" when X = 13 AND Y = 0 else
"1111111100000" when X = 14 AND Y = 0 else
"1111111100000" when X = 15 AND Y = 0 else
"1111111100000" when X = 16 AND Y = 0 else
"1111111100000" when X = 17 AND Y = 0 else
"1111111100000" when X = 18 AND Y = 0 else
"1111111100000" when X = 19 AND Y = 0 else
"1111111100000" when X = 20 AND Y = 0 else
"1111111100000" when X = 21 AND Y = 0 else
"1111111100000" when X = 22 AND Y = 0 else
"1111111100000" when X = 23 AND Y = 0 else
"1111111100000" when X = 24 AND Y = 0 else
"1111111100000" when X = 25 AND Y = 0 else
"1111111100000" when X = 26 AND Y = 0 else
"1111111100000" when X = 27 AND Y = 0 else
"1111111100000" when X = 28 AND Y = 0 else
"1111111100000" when X = 29 AND Y = 0 else
"1111111100000" when X = 30 AND Y = 0 else
"1111111100000" when X = 31 AND Y = 0 else
"1111111100000" when X = 32 AND Y = 0 else
"1111111100000" when X = 33 AND Y = 0 else
"1111111100000" when X = 34 AND Y = 0 else
"1111111100000" when X = 35 AND Y = 0 else
"1111111100000" when X = 36 AND Y = 0 else
"1111111100000" when X = 37 AND Y = 0 else
"1111111100000" when X = 38 AND Y = 0 else
"1111111100000" when X = 39 AND Y = 0 else
"1111111100000" when X = 40 AND Y = 0 else
"1111111100000" when X = 41 AND Y = 0 else
"1111111100000" when X = 42 AND Y = 0 else
"1111111100000" when X = 43 AND Y = 0 else
"1111111100000" when X = 44 AND Y = 0 else
"1111111100000" when X = 45 AND Y = 0 else
"1111111100000" when X = 0 AND Y = 1 else
"1111111100000" when X = 1 AND Y = 1 else
"1111111100000" when X = 2 AND Y = 1 else
"1111111100000" when X = 3 AND Y = 1 else
"1111111100000" when X = 4 AND Y = 1 else
"1111111100000" when X = 5 AND Y = 1 else
"1111111100000" when X = 6 AND Y = 1 else
"1111111100000" when X = 7 AND Y = 1 else
"1111111100000" when X = 8 AND Y = 1 else
"1111111100000" when X = 9 AND Y = 1 else
"1111111100000" when X = 10 AND Y = 1 else
"1111111100000" when X = 11 AND Y = 1 else
"1111111100000" when X = 12 AND Y = 1 else
"1111111100000" when X = 13 AND Y = 1 else
"1111111100000" when X = 14 AND Y = 1 else
"1111111100000" when X = 15 AND Y = 1 else
"1111111100000" when X = 16 AND Y = 1 else
"1111111100000" when X = 17 AND Y = 1 else
"1111111100000" when X = 18 AND Y = 1 else
"1111111100000" when X = 19 AND Y = 1 else
"1111111100000" when X = 20 AND Y = 1 else
"1111111100000" when X = 21 AND Y = 1 else
"1111111100000" when X = 22 AND Y = 1 else
"1111111100000" when X = 23 AND Y = 1 else
"1111111100000" when X = 24 AND Y = 1 else
"1111111100000" when X = 25 AND Y = 1 else
"1111111100000" when X = 26 AND Y = 1 else
"1111111100000" when X = 27 AND Y = 1 else
"1111111100000" when X = 28 AND Y = 1 else
"1111111100000" when X = 29 AND Y = 1 else
"1111111100000" when X = 30 AND Y = 1 else
"1111111100000" when X = 31 AND Y = 1 else
"1111111100000" when X = 32 AND Y = 1 else
"1111111100000" when X = 33 AND Y = 1 else
"1111111100000" when X = 34 AND Y = 1 else
"1111111100000" when X = 35 AND Y = 1 else
"1111111100000" when X = 36 AND Y = 1 else
"1111111100000" when X = 37 AND Y = 1 else
"1111111100000" when X = 38 AND Y = 1 else
"1111111100000" when X = 39 AND Y = 1 else
"1111111100000" when X = 40 AND Y = 1 else
"1111111100000" when X = 41 AND Y = 1 else
"1111111100000" when X = 42 AND Y = 1 else
"1111111100000" when X = 43 AND Y = 1 else
"1111111100000" when X = 44 AND Y = 1 else
"1111111100000" when X = 45 AND Y = 1 else
"1111111100000" when X = 0 AND Y = 2 else
"1111111100000" when X = 1 AND Y = 2 else
"1111111100000" when X = 2 AND Y = 2 else
"1111111100000" when X = 3 AND Y = 2 else
"1111111100000" when X = 4 AND Y = 2 else
"1111111100000" when X = 5 AND Y = 2 else
"1111111100000" when X = 6 AND Y = 2 else
"1111111100000" when X = 7 AND Y = 2 else
"1111111100000" when X = 8 AND Y = 2 else
"1111111100000" when X = 9 AND Y = 2 else
"1111111100000" when X = 10 AND Y = 2 else
"1111111100000" when X = 11 AND Y = 2 else
"1111111100000" when X = 12 AND Y = 2 else
"1111111100000" when X = 13 AND Y = 2 else
"1111111100000" when X = 14 AND Y = 2 else
"1111111100000" when X = 15 AND Y = 2 else
"1111111100000" when X = 16 AND Y = 2 else
"1111111100000" when X = 17 AND Y = 2 else
"1111111100000" when X = 18 AND Y = 2 else
"1111111100000" when X = 19 AND Y = 2 else
"1111111100000" when X = 20 AND Y = 2 else
"1111111100000" when X = 21 AND Y = 2 else
"1111111100000" when X = 22 AND Y = 2 else
"1111111100000" when X = 23 AND Y = 2 else
"1111111100000" when X = 24 AND Y = 2 else
"1111111100000" when X = 25 AND Y = 2 else
"1111111100000" when X = 26 AND Y = 2 else
"1111111100000" when X = 27 AND Y = 2 else
"1111111100000" when X = 28 AND Y = 2 else
"1111111100000" when X = 29 AND Y = 2 else
"1111111100000" when X = 30 AND Y = 2 else
"1111111100000" when X = 31 AND Y = 2 else
"1111111100000" when X = 32 AND Y = 2 else
"1111111100000" when X = 33 AND Y = 2 else
"1111111100000" when X = 34 AND Y = 2 else
"1111111100000" when X = 35 AND Y = 2 else
"1111111100000" when X = 36 AND Y = 2 else
"1111111100000" when X = 37 AND Y = 2 else
"1111111100000" when X = 38 AND Y = 2 else
"1111111100000" when X = 39 AND Y = 2 else
"1111111100000" when X = 40 AND Y = 2 else
"1111111100000" when X = 41 AND Y = 2 else
"1111111100000" when X = 42 AND Y = 2 else
"1111111100000" when X = 43 AND Y = 2 else
"1111111100000" when X = 44 AND Y = 2 else
"1111111100000" when X = 45 AND Y = 2 else
"1111111100000" when X = 0 AND Y = 3 else
"1111111100000" when X = 1 AND Y = 3 else
"1111111100000" when X = 2 AND Y = 3 else
"1111111100000" when X = 3 AND Y = 3 else
"1111111100000" when X = 4 AND Y = 3 else
"1111111100000" when X = 5 AND Y = 3 else
"1111111100000" when X = 6 AND Y = 3 else
"1111111100000" when X = 7 AND Y = 3 else
"1111111100000" when X = 8 AND Y = 3 else
"1111111100000" when X = 9 AND Y = 3 else
"1111111100000" when X = 10 AND Y = 3 else
"1111111100000" when X = 11 AND Y = 3 else
"1111111100000" when X = 12 AND Y = 3 else
"1111111100000" when X = 13 AND Y = 3 else
"1111111100000" when X = 14 AND Y = 3 else
"1111111100000" when X = 15 AND Y = 3 else
"1111111100000" when X = 16 AND Y = 3 else
"1111111100000" when X = 17 AND Y = 3 else
"1111111100000" when X = 18 AND Y = 3 else
"1111111100000" when X = 19 AND Y = 3 else
"0111101111101" when X = 20 AND Y = 3 else
"0100011011111" when X = 21 AND Y = 3 else
"0100011011111" when X = 22 AND Y = 3 else
"0100011111111" when X = 23 AND Y = 3 else
"1111111100001" when X = 24 AND Y = 3 else
"1111111100000" when X = 25 AND Y = 3 else
"1111111100000" when X = 26 AND Y = 3 else
"1111111100000" when X = 27 AND Y = 3 else
"1111111100000" when X = 28 AND Y = 3 else
"1111111100000" when X = 29 AND Y = 3 else
"1111111100000" when X = 30 AND Y = 3 else
"1111111100000" when X = 31 AND Y = 3 else
"1111111100000" when X = 32 AND Y = 3 else
"1111111100000" when X = 33 AND Y = 3 else
"1111111100000" when X = 34 AND Y = 3 else
"1111111100000" when X = 35 AND Y = 3 else
"1111111100000" when X = 36 AND Y = 3 else
"1111111100000" when X = 37 AND Y = 3 else
"1111111100000" when X = 38 AND Y = 3 else
"1111111100000" when X = 39 AND Y = 3 else
"1111111100000" when X = 40 AND Y = 3 else
"1111111100000" when X = 41 AND Y = 3 else
"1111111100000" when X = 42 AND Y = 3 else
"1111111100000" when X = 43 AND Y = 3 else
"1111111100000" when X = 44 AND Y = 3 else
"1111111100000" when X = 45 AND Y = 3 else
"1111111100000" when X = 0 AND Y = 4 else
"1111111100000" when X = 1 AND Y = 4 else
"1111111100000" when X = 2 AND Y = 4 else
"1111111100000" when X = 3 AND Y = 4 else
"1111111100000" when X = 4 AND Y = 4 else
"1111111100000" when X = 5 AND Y = 4 else
"1111111100000" when X = 6 AND Y = 4 else
"1111111100000" when X = 7 AND Y = 4 else
"1111111100000" when X = 8 AND Y = 4 else
"1111111100000" when X = 9 AND Y = 4 else
"1111111100000" when X = 10 AND Y = 4 else
"1111111100000" when X = 11 AND Y = 4 else
"1111111100000" when X = 12 AND Y = 4 else
"1111111100000" when X = 13 AND Y = 4 else
"1111111100000" when X = 14 AND Y = 4 else
"1111111100000" when X = 15 AND Y = 4 else
"1111111100000" when X = 16 AND Y = 4 else
"1111111100000" when X = 17 AND Y = 4 else
"1111111100000" when X = 18 AND Y = 4 else
"1000101111101" when X = 19 AND Y = 4 else
"0010010111111" when X = 20 AND Y = 4 else
"0010010111111" when X = 21 AND Y = 4 else
"0101101011111" when X = 22 AND Y = 4 else
"0001010011111" when X = 23 AND Y = 4 else
"0011011011111" when X = 24 AND Y = 4 else
"1111111100001" when X = 25 AND Y = 4 else
"1111111100000" when X = 26 AND Y = 4 else
"1111111100000" when X = 27 AND Y = 4 else
"1111111100000" when X = 28 AND Y = 4 else
"1111111100000" when X = 29 AND Y = 4 else
"1111111100000" when X = 30 AND Y = 4 else
"1111111100000" when X = 31 AND Y = 4 else
"1111111100000" when X = 32 AND Y = 4 else
"1111111100000" when X = 33 AND Y = 4 else
"1111111100000" when X = 34 AND Y = 4 else
"1111111100000" when X = 35 AND Y = 4 else
"1111111100000" when X = 36 AND Y = 4 else
"1111111100000" when X = 37 AND Y = 4 else
"1111111100000" when X = 38 AND Y = 4 else
"1111111100000" when X = 39 AND Y = 4 else
"1111111100000" when X = 40 AND Y = 4 else
"1111111100000" when X = 41 AND Y = 4 else
"1111111100000" when X = 42 AND Y = 4 else
"1111111100000" when X = 43 AND Y = 4 else
"1111111100000" when X = 44 AND Y = 4 else
"1111111100000" when X = 45 AND Y = 4 else
"1111111100000" when X = 0 AND Y = 5 else
"1111111100000" when X = 1 AND Y = 5 else
"1111111100000" when X = 2 AND Y = 5 else
"1111111100000" when X = 3 AND Y = 5 else
"1111111100000" when X = 4 AND Y = 5 else
"1111111100000" when X = 5 AND Y = 5 else
"1111111100000" when X = 6 AND Y = 5 else
"0111101010111" when X = 7 AND Y = 5 else
"0111101010101" when X = 8 AND Y = 5 else
"0111101010111" when X = 9 AND Y = 5 else
"1000110011001" when X = 10 AND Y = 5 else
"1111111100000" when X = 11 AND Y = 5 else
"1111111100000" when X = 12 AND Y = 5 else
"1111111100000" when X = 13 AND Y = 5 else
"1111111100000" when X = 14 AND Y = 5 else
"1111111100000" when X = 15 AND Y = 5 else
"1011110011001" when X = 16 AND Y = 5 else
"1011101110111" when X = 17 AND Y = 5 else
"1001110011011" when X = 18 AND Y = 5 else
"0010010111111" when X = 19 AND Y = 5 else
"0001001111101" when X = 20 AND Y = 5 else
"0110110010111" when X = 21 AND Y = 5 else
"0111110110101" when X = 22 AND Y = 5 else
"0101101110111" when X = 23 AND Y = 5 else
"0001001011111" when X = 24 AND Y = 5 else
"0011011111111" when X = 25 AND Y = 5 else
"1010110011001" when X = 26 AND Y = 5 else
"1011101110111" when X = 27 AND Y = 5 else
"1011110011001" when X = 28 AND Y = 5 else
"1111111100000" when X = 29 AND Y = 5 else
"1111111100000" when X = 30 AND Y = 5 else
"1111111100000" when X = 31 AND Y = 5 else
"1111111100000" when X = 32 AND Y = 5 else
"1111111100000" when X = 33 AND Y = 5 else
"1000110011001" when X = 34 AND Y = 5 else
"0111101010101" when X = 35 AND Y = 5 else
"0111101010101" when X = 36 AND Y = 5 else
"0111101111001" when X = 37 AND Y = 5 else
"1111111100000" when X = 38 AND Y = 5 else
"1111111100000" when X = 39 AND Y = 5 else
"1111111100000" when X = 40 AND Y = 5 else
"1111111100000" when X = 41 AND Y = 5 else
"1111111100000" when X = 42 AND Y = 5 else
"1111111100000" when X = 43 AND Y = 5 else
"1111111100000" when X = 44 AND Y = 5 else
"1111111100000" when X = 45 AND Y = 5 else
"1111111100000" when X = 0 AND Y = 6 else
"1111111100000" when X = 1 AND Y = 6 else
"1111111100000" when X = 2 AND Y = 6 else
"1111111100000" when X = 3 AND Y = 6 else
"1111111100000" when X = 4 AND Y = 6 else
"1111111100000" when X = 5 AND Y = 6 else
"0111100110101" when X = 6 AND Y = 6 else
"0100010101011" when X = 7 AND Y = 6 else
"0011001100111" when X = 8 AND Y = 6 else
"0000000000001" when X = 9 AND Y = 6 else
"0010010001001" when X = 10 AND Y = 6 else
"1000101111001" when X = 11 AND Y = 6 else
"1111111100000" when X = 12 AND Y = 6 else
"1000100111001" when X = 13 AND Y = 6 else
"1000100011001" when X = 14 AND Y = 6 else
"1011101010101" when X = 15 AND Y = 6 else
"1111100100111" when X = 16 AND Y = 6 else
"1111010000011" when X = 17 AND Y = 6 else
"1010100010001" when X = 18 AND Y = 6 else
"0000010011111" when X = 19 AND Y = 6 else
"0011010011011" when X = 20 AND Y = 6 else
"1110111000111" when X = 21 AND Y = 6 else
"1110111100011" when X = 22 AND Y = 6 else
"1100110101011" when X = 23 AND Y = 6 else
"0001001011101" when X = 24 AND Y = 6 else
"0000011011101" when X = 25 AND Y = 6 else
"1100011101101" when X = 26 AND Y = 6 else
"1111010000001" when X = 27 AND Y = 6 else
"1111100100111" when X = 28 AND Y = 6 else
"1011101010101" when X = 29 AND Y = 6 else
"1000100011001" when X = 30 AND Y = 6 else
"1000100111001" when X = 31 AND Y = 6 else
"1111111100000" when X = 32 AND Y = 6 else
"1000110011001" when X = 33 AND Y = 6 else
"0011010001001" when X = 34 AND Y = 6 else
"0000000000001" when X = 35 AND Y = 6 else
"0011001100111" when X = 36 AND Y = 6 else
"0100010101011" when X = 37 AND Y = 6 else
"0111101010111" when X = 38 AND Y = 6 else
"1111111100000" when X = 39 AND Y = 6 else
"1111111100000" when X = 40 AND Y = 6 else
"1111111100000" when X = 41 AND Y = 6 else
"1111111100000" when X = 42 AND Y = 6 else
"1111111100000" when X = 43 AND Y = 6 else
"1111111100000" when X = 44 AND Y = 6 else
"1111111100000" when X = 45 AND Y = 6 else
"1111111100000" when X = 0 AND Y = 7 else
"1111111100000" when X = 1 AND Y = 7 else
"1111111100000" when X = 2 AND Y = 7 else
"1111111100000" when X = 3 AND Y = 7 else
"1111111100000" when X = 4 AND Y = 7 else
"1111111100000" when X = 5 AND Y = 7 else
"0011010101011" when X = 6 AND Y = 7 else
"0011001100111" when X = 7 AND Y = 7 else
"0010001000101" when X = 8 AND Y = 7 else
"0000000000001" when X = 9 AND Y = 7 else
"0000000000001" when X = 10 AND Y = 7 else
"0101010001111" when X = 11 AND Y = 7 else
"1000010110111" when X = 12 AND Y = 7 else
"1001001110001" when X = 13 AND Y = 7 else
"1100010101011" when X = 14 AND Y = 7 else
"1110100000101" when X = 15 AND Y = 7 else
"1111011100001" when X = 16 AND Y = 7 else
"1101010001001" when X = 17 AND Y = 7 else
"0101011111001" when X = 18 AND Y = 7 else
"0001001111111" when X = 19 AND Y = 7 else
"1000100110011" when X = 20 AND Y = 7 else
"1110111000011" when X = 21 AND Y = 7 else
"1111111100001" when X = 22 AND Y = 7 else
"1110111000101" when X = 23 AND Y = 7 else
"0111100010101" when X = 24 AND Y = 7 else
"0001001111111" when X = 25 AND Y = 7 else
"0110100010111" when X = 26 AND Y = 7 else
"1101010101001" when X = 27 AND Y = 7 else
"1111011100001" when X = 28 AND Y = 7 else
"1110100000101" when X = 29 AND Y = 7 else
"1100010101011" when X = 30 AND Y = 7 else
"1001001110001" when X = 31 AND Y = 7 else
"1000010110111" when X = 32 AND Y = 7 else
"0110010001111" when X = 33 AND Y = 7 else
"0000000000001" when X = 34 AND Y = 7 else
"0000000000001" when X = 35 AND Y = 7 else
"0011001100111" when X = 36 AND Y = 7 else
"0010001000101" when X = 37 AND Y = 7 else
"0101011101111" when X = 38 AND Y = 7 else
"1111111100000" when X = 39 AND Y = 7 else
"1111111100000" when X = 40 AND Y = 7 else
"1111111100000" when X = 41 AND Y = 7 else
"1111111100000" when X = 42 AND Y = 7 else
"1111111100000" when X = 43 AND Y = 7 else
"1111111100000" when X = 44 AND Y = 7 else
"1111111100000" when X = 45 AND Y = 7 else
"1111111100000" when X = 0 AND Y = 8 else
"1111111100000" when X = 1 AND Y = 8 else
"1111111100000" when X = 2 AND Y = 8 else
"1111111100000" when X = 3 AND Y = 8 else
"1111111100000" when X = 4 AND Y = 8 else
"1111111100000" when X = 5 AND Y = 8 else
"0011010101011" when X = 6 AND Y = 8 else
"0000000000001" when X = 7 AND Y = 8 else
"0000000000001" when X = 8 AND Y = 8 else
"0000000000001" when X = 9 AND Y = 8 else
"0110001100001" when X = 10 AND Y = 8 else
"1101011100111" when X = 11 AND Y = 8 else
"1101011001001" when X = 12 AND Y = 8 else
"1110011100111" when X = 13 AND Y = 8 else
"1111100100001" when X = 14 AND Y = 8 else
"1111100100001" when X = 15 AND Y = 8 else
"1111011100001" when X = 16 AND Y = 8 else
"1011011101101" when X = 17 AND Y = 8 else
"0000011011111" when X = 18 AND Y = 8 else
"0010001111011" when X = 19 AND Y = 8 else
"1101110101001" when X = 20 AND Y = 8 else
"1111111000001" when X = 21 AND Y = 8 else
"1111111000001" when X = 22 AND Y = 8 else
"1111111000001" when X = 23 AND Y = 8 else
"1011101101101" when X = 24 AND Y = 8 else
"0001000111101" when X = 25 AND Y = 8 else
"0000100011101" when X = 26 AND Y = 8 else
"1011100001101" when X = 27 AND Y = 8 else
"1111011100001" when X = 28 AND Y = 8 else
"1111100100001" when X = 29 AND Y = 8 else
"1111100100001" when X = 30 AND Y = 8 else
"1110011100111" when X = 31 AND Y = 8 else
"1101011001001" when X = 32 AND Y = 8 else
"1101011100111" when X = 33 AND Y = 8 else
"0110001100001" when X = 34 AND Y = 8 else
"0000000000001" when X = 35 AND Y = 8 else
"0000000000001" when X = 36 AND Y = 8 else
"0000000000001" when X = 37 AND Y = 8 else
"0101011101111" when X = 38 AND Y = 8 else
"1111111100000" when X = 39 AND Y = 8 else
"1111111100000" when X = 40 AND Y = 8 else
"1111111100000" when X = 41 AND Y = 8 else
"1111111100000" when X = 42 AND Y = 8 else
"1111111100000" when X = 43 AND Y = 8 else
"1111111100000" when X = 44 AND Y = 8 else
"1111111100000" when X = 45 AND Y = 8 else
"1111111100000" when X = 0 AND Y = 9 else
"1111111100000" when X = 1 AND Y = 9 else
"1111111100000" when X = 2 AND Y = 9 else
"1111111100000" when X = 3 AND Y = 9 else
"1111111100000" when X = 4 AND Y = 9 else
"1111111100000" when X = 5 AND Y = 9 else
"0011010101011" when X = 6 AND Y = 9 else
"0000000000001" when X = 7 AND Y = 9 else
"0001000000001" when X = 8 AND Y = 9 else
"0111001100001" when X = 9 AND Y = 9 else
"1110100000001" when X = 10 AND Y = 9 else
"1111100000001" when X = 11 AND Y = 9 else
"1111100000001" when X = 12 AND Y = 9 else
"1111100100001" when X = 13 AND Y = 9 else
"1111100100001" when X = 14 AND Y = 9 else
"1111100100001" when X = 15 AND Y = 9 else
"1101100101001" when X = 16 AND Y = 9 else
"0100110011001" when X = 17 AND Y = 9 else
"0011100011001" when X = 18 AND Y = 9 else
"1011011101101" when X = 19 AND Y = 9 else
"1111100100001" when X = 20 AND Y = 9 else
"1111100100001" when X = 21 AND Y = 9 else
"1111100100001" when X = 22 AND Y = 9 else
"1111100100001" when X = 23 AND Y = 9 else
"1111100100011" when X = 24 AND Y = 9 else
"1001011010001" when X = 25 AND Y = 9 else
"0010100111011" when X = 26 AND Y = 9 else
"0100110011001" when X = 27 AND Y = 9 else
"1101100101001" when X = 28 AND Y = 9 else
"1111100100001" when X = 29 AND Y = 9 else
"1111100100001" when X = 30 AND Y = 9 else
"1111100100001" when X = 31 AND Y = 9 else
"1111100000001" when X = 32 AND Y = 9 else
"1111100000001" when X = 33 AND Y = 9 else
"1111100000001" when X = 34 AND Y = 9 else
"0110001100001" when X = 35 AND Y = 9 else
"0000000000001" when X = 36 AND Y = 9 else
"0000000000001" when X = 37 AND Y = 9 else
"0101011101111" when X = 38 AND Y = 9 else
"1111111100000" when X = 39 AND Y = 9 else
"1111111100000" when X = 40 AND Y = 9 else
"1111111100000" when X = 41 AND Y = 9 else
"1111111100000" when X = 42 AND Y = 9 else
"1111111100000" when X = 43 AND Y = 9 else
"1111111100000" when X = 44 AND Y = 9 else
"1111111100000" when X = 45 AND Y = 9 else
"1111111100000" when X = 0 AND Y = 10 else
"1111111100000" when X = 1 AND Y = 10 else
"1111111100000" when X = 2 AND Y = 10 else
"1111111100000" when X = 3 AND Y = 10 else
"1111111100000" when X = 4 AND Y = 10 else
"1111111100000" when X = 5 AND Y = 10 else
"0011010001011" when X = 6 AND Y = 10 else
"0000000000001" when X = 7 AND Y = 10 else
"1000010000001" when X = 8 AND Y = 10 else
"1111100000001" when X = 9 AND Y = 10 else
"1111100000001" when X = 10 AND Y = 10 else
"1111010000001" when X = 11 AND Y = 10 else
"1111010100001" when X = 12 AND Y = 10 else
"1111011000001" when X = 13 AND Y = 10 else
"1111011000001" when X = 14 AND Y = 10 else
"1111011000001" when X = 15 AND Y = 10 else
"1110011000111" when X = 16 AND Y = 10 else
"1001100010001" when X = 17 AND Y = 10 else
"1101011101011" when X = 18 AND Y = 10 else
"1111011000001" when X = 19 AND Y = 10 else
"1111011000001" when X = 20 AND Y = 10 else
"1111011000001" when X = 21 AND Y = 10 else
"1111011000001" when X = 22 AND Y = 10 else
"1111011000001" when X = 23 AND Y = 10 else
"1111011000001" when X = 24 AND Y = 10 else
"1111011000001" when X = 25 AND Y = 10 else
"1011011101101" when X = 26 AND Y = 10 else
"1001100010001" when X = 27 AND Y = 10 else
"1110011000111" when X = 28 AND Y = 10 else
"1111011000001" when X = 29 AND Y = 10 else
"1111011000001" when X = 30 AND Y = 10 else
"1111011000001" when X = 31 AND Y = 10 else
"1111010100001" when X = 32 AND Y = 10 else
"1111010000001" when X = 33 AND Y = 10 else
"1111100000001" when X = 34 AND Y = 10 else
"1111100000001" when X = 35 AND Y = 10 else
"0110001100001" when X = 36 AND Y = 10 else
"0000000000001" when X = 37 AND Y = 10 else
"0101011101111" when X = 38 AND Y = 10 else
"1111111100000" when X = 39 AND Y = 10 else
"1111111100000" when X = 40 AND Y = 10 else
"1111111100000" when X = 41 AND Y = 10 else
"1111111100000" when X = 42 AND Y = 10 else
"1111111100000" when X = 43 AND Y = 10 else
"1111111100000" when X = 44 AND Y = 10 else
"1111111100000" when X = 45 AND Y = 10 else
"1111111100000" when X = 0 AND Y = 11 else
"1111111100000" when X = 1 AND Y = 11 else
"1111111100000" when X = 2 AND Y = 11 else
"1111111100000" when X = 3 AND Y = 11 else
"1111111100000" when X = 4 AND Y = 11 else
"1011110010111" when X = 5 AND Y = 11 else
"1010011000111" when X = 6 AND Y = 11 else
"1001010100001" when X = 7 AND Y = 11 else
"1110100000001" when X = 8 AND Y = 11 else
"1111100000001" when X = 9 AND Y = 11 else
"1111100000001" when X = 10 AND Y = 11 else
"1111010000001" when X = 11 AND Y = 11 else
"1100000000001" when X = 12 AND Y = 11 else
"1011000000001" when X = 13 AND Y = 11 else
"1011000000001" when X = 14 AND Y = 11 else
"1011000000001" when X = 15 AND Y = 11 else
"1011000000001" when X = 16 AND Y = 11 else
"1011000000001" when X = 17 AND Y = 11 else
"1011000000001" when X = 18 AND Y = 11 else
"1011000000001" when X = 19 AND Y = 11 else
"1011000000001" when X = 20 AND Y = 11 else
"1011000000001" when X = 21 AND Y = 11 else
"1011000000001" when X = 22 AND Y = 11 else
"1011000000001" when X = 23 AND Y = 11 else
"1011000000001" when X = 24 AND Y = 11 else
"1011000000001" when X = 25 AND Y = 11 else
"1011000000001" when X = 26 AND Y = 11 else
"1011000000001" when X = 27 AND Y = 11 else
"1011000000001" when X = 28 AND Y = 11 else
"1011000000001" when X = 29 AND Y = 11 else
"1011000000001" when X = 30 AND Y = 11 else
"1011000000001" when X = 31 AND Y = 11 else
"1100000000001" when X = 32 AND Y = 11 else
"1111010000001" when X = 33 AND Y = 11 else
"1111100000001" when X = 34 AND Y = 11 else
"1111100000001" when X = 35 AND Y = 11 else
"1110100000001" when X = 36 AND Y = 11 else
"1001010100001" when X = 37 AND Y = 11 else
"1011100001001" when X = 38 AND Y = 11 else
"1010110011001" when X = 39 AND Y = 11 else
"1111111100000" when X = 40 AND Y = 11 else
"1111111100000" when X = 41 AND Y = 11 else
"1111111100000" when X = 42 AND Y = 11 else
"1111111100000" when X = 43 AND Y = 11 else
"1111111100000" when X = 44 AND Y = 11 else
"1111111100000" when X = 45 AND Y = 11 else
"1111111100000" when X = 0 AND Y = 12 else
"1111111100000" when X = 1 AND Y = 12 else
"0101011101111" when X = 2 AND Y = 12 else
"0010001100111" when X = 3 AND Y = 12 else
"0010001100111" when X = 4 AND Y = 12 else
"0011001000101" when X = 5 AND Y = 12 else
"0100001000001" when X = 6 AND Y = 12 else
"0100001000001" when X = 7 AND Y = 12 else
"0011001000001" when X = 8 AND Y = 12 else
"0111010000001" when X = 9 AND Y = 12 else
"1111100000001" when X = 10 AND Y = 12 else
"1111010000001" when X = 11 AND Y = 12 else
"1010000000001" when X = 12 AND Y = 12 else
"1000000000001" when X = 13 AND Y = 12 else
"1000000000001" when X = 14 AND Y = 12 else
"1000000000001" when X = 15 AND Y = 12 else
"1000000000001" when X = 16 AND Y = 12 else
"1000000000001" when X = 17 AND Y = 12 else
"1000000000001" when X = 18 AND Y = 12 else
"1000000000001" when X = 19 AND Y = 12 else
"1000000000001" when X = 20 AND Y = 12 else
"1000000000001" when X = 21 AND Y = 12 else
"1001000000001" when X = 22 AND Y = 12 else
"1000000000001" when X = 23 AND Y = 12 else
"1000000000001" when X = 24 AND Y = 12 else
"1000000000001" when X = 25 AND Y = 12 else
"1000000000001" when X = 26 AND Y = 12 else
"1000000000001" when X = 27 AND Y = 12 else
"1000000000001" when X = 28 AND Y = 12 else
"1000000000001" when X = 29 AND Y = 12 else
"1000000000001" when X = 30 AND Y = 12 else
"1000000000001" when X = 31 AND Y = 12 else
"1010000000001" when X = 32 AND Y = 12 else
"1111010000001" when X = 33 AND Y = 12 else
"1111100000001" when X = 34 AND Y = 12 else
"0111010000001" when X = 35 AND Y = 12 else
"0011001000001" when X = 36 AND Y = 12 else
"0100001000001" when X = 37 AND Y = 12 else
"0100001000001" when X = 38 AND Y = 12 else
"0010001100101" when X = 39 AND Y = 12 else
"0010001100111" when X = 40 AND Y = 12 else
"0010001100111" when X = 41 AND Y = 12 else
"0110100010011" when X = 42 AND Y = 12 else
"1111111100000" when X = 43 AND Y = 12 else
"1111111100000" when X = 44 AND Y = 12 else
"1111111100000" when X = 45 AND Y = 12 else
"1111111100000" when X = 0 AND Y = 13 else
"0110100110101" when X = 1 AND Y = 13 else
"0000000100011" when X = 2 AND Y = 13 else
"0000000000001" when X = 3 AND Y = 13 else
"0000000000001" when X = 4 AND Y = 13 else
"0000000000001" when X = 5 AND Y = 13 else
"0001000100011" when X = 6 AND Y = 13 else
"0001000100011" when X = 7 AND Y = 13 else
"0000000000001" when X = 8 AND Y = 13 else
"0001000000001" when X = 9 AND Y = 13 else
"1000010100101" when X = 10 AND Y = 13 else
"1111001100011" when X = 11 AND Y = 13 else
"1010000000001" when X = 12 AND Y = 13 else
"1001000000001" when X = 13 AND Y = 13 else
"1001000000001" when X = 14 AND Y = 13 else
"1001000000001" when X = 15 AND Y = 13 else
"1001000000001" when X = 16 AND Y = 13 else
"1001000000001" when X = 17 AND Y = 13 else
"1001000000001" when X = 18 AND Y = 13 else
"1001000000001" when X = 19 AND Y = 13 else
"1000000000001" when X = 20 AND Y = 13 else
"1011000000001" when X = 21 AND Y = 13 else
"1110000000001" when X = 22 AND Y = 13 else
"1010000000001" when X = 23 AND Y = 13 else
"1000000000001" when X = 24 AND Y = 13 else
"1001000000001" when X = 25 AND Y = 13 else
"1001000000001" when X = 26 AND Y = 13 else
"1001000000001" when X = 27 AND Y = 13 else
"1001000000001" when X = 28 AND Y = 13 else
"1001000000001" when X = 29 AND Y = 13 else
"1001000000001" when X = 30 AND Y = 13 else
"1001000000001" when X = 31 AND Y = 13 else
"1010000000001" when X = 32 AND Y = 13 else
"1111001100011" when X = 33 AND Y = 13 else
"1001010100101" when X = 34 AND Y = 13 else
"0001000000001" when X = 35 AND Y = 13 else
"0000000000011" when X = 36 AND Y = 13 else
"0001000100011" when X = 37 AND Y = 13 else
"0001000100011" when X = 38 AND Y = 13 else
"0000000000001" when X = 39 AND Y = 13 else
"0001000000001" when X = 40 AND Y = 13 else
"0000000000001" when X = 41 AND Y = 13 else
"0001001000101" when X = 42 AND Y = 13 else
"0111101010111" when X = 43 AND Y = 13 else
"1111111100000" when X = 44 AND Y = 13 else
"1111111100000" when X = 45 AND Y = 13 else
"1111111100000" when X = 0 AND Y = 14 else
"0101011110001" when X = 1 AND Y = 14 else
"0000000000001" when X = 2 AND Y = 14 else
"0100010001001" when X = 3 AND Y = 14 else
"0100010001001" when X = 4 AND Y = 14 else
"0010001000101" when X = 5 AND Y = 14 else
"0110011001101" when X = 6 AND Y = 14 else
"0110011001101" when X = 7 AND Y = 14 else
"0100010001001" when X = 8 AND Y = 14 else
"0000000000001" when X = 9 AND Y = 14 else
"0001000101111" when X = 10 AND Y = 14 else
"1010001001101" when X = 11 AND Y = 14 else
"1000000100111" when X = 12 AND Y = 14 else
"0110000001001" when X = 13 AND Y = 14 else
"0110000001001" when X = 14 AND Y = 14 else
"0110000001001" when X = 15 AND Y = 14 else
"0110000001001" when X = 16 AND Y = 14 else
"0110000001001" when X = 17 AND Y = 14 else
"0110000001001" when X = 18 AND Y = 14 else
"0110000001001" when X = 19 AND Y = 14 else
"0111000000111" when X = 20 AND Y = 14 else
"1100000000001" when X = 21 AND Y = 14 else
"1111000000001" when X = 22 AND Y = 14 else
"1011000000011" when X = 23 AND Y = 14 else
"0110000001001" when X = 24 AND Y = 14 else
"0110000001001" when X = 25 AND Y = 14 else
"0110000001001" when X = 26 AND Y = 14 else
"0110000001001" when X = 27 AND Y = 14 else
"0110000001001" when X = 28 AND Y = 14 else
"0110000001001" when X = 29 AND Y = 14 else
"0110000001001" when X = 30 AND Y = 14 else
"0110000001001" when X = 31 AND Y = 14 else
"1000000100111" when X = 32 AND Y = 14 else
"1010001001101" when X = 33 AND Y = 14 else
"0001000101111" when X = 34 AND Y = 14 else
"0000000000001" when X = 35 AND Y = 14 else
"0101010101011" when X = 36 AND Y = 14 else
"0110011001101" when X = 37 AND Y = 14 else
"0110011001101" when X = 38 AND Y = 14 else
"0010001000101" when X = 39 AND Y = 14 else
"0101010101011" when X = 40 AND Y = 14 else
"0011001100111" when X = 41 AND Y = 14 else
"0000000000001" when X = 42 AND Y = 14 else
"0111101010101" when X = 43 AND Y = 14 else
"1111111100000" when X = 44 AND Y = 14 else
"1111111100000" when X = 45 AND Y = 14 else
"1111111100000" when X = 0 AND Y = 15 else
"0101011110001" when X = 1 AND Y = 15 else
"0000000000001" when X = 2 AND Y = 15 else
"0000000000001" when X = 3 AND Y = 15 else
"0000000000001" when X = 4 AND Y = 15 else
"0000000000001" when X = 5 AND Y = 15 else
"0000000000001" when X = 6 AND Y = 15 else
"0000000000001" when X = 7 AND Y = 15 else
"0000000000001" when X = 8 AND Y = 15 else
"0000000000001" when X = 9 AND Y = 15 else
"0000000001111" when X = 10 AND Y = 15 else
"1001000101111" when X = 11 AND Y = 15 else
"0011000111001" when X = 12 AND Y = 15 else
"0001001011101" when X = 13 AND Y = 15 else
"0000010011001" when X = 14 AND Y = 15 else
"0000010011001" when X = 15 AND Y = 15 else
"0001010011001" when X = 16 AND Y = 15 else
"0011000111001" when X = 17 AND Y = 15 else
"0010001111001" when X = 18 AND Y = 15 else
"0010001011011" when X = 19 AND Y = 15 else
"0110000110101" when X = 20 AND Y = 15 else
"1111000000011" when X = 21 AND Y = 15 else
"1111000000001" when X = 22 AND Y = 15 else
"1110000000101" when X = 23 AND Y = 15 else
"0100000110111" when X = 24 AND Y = 15 else
"0010001011001" when X = 25 AND Y = 15 else
"0010001011001" when X = 26 AND Y = 15 else
"0011000111001" when X = 27 AND Y = 15 else
"0001010011001" when X = 28 AND Y = 15 else
"0000010011001" when X = 29 AND Y = 15 else
"0001010011001" when X = 30 AND Y = 15 else
"0001001011101" when X = 31 AND Y = 15 else
"0011000111011" when X = 32 AND Y = 15 else
"1001000101111" when X = 33 AND Y = 15 else
"0000000001111" when X = 34 AND Y = 15 else
"0000000000001" when X = 35 AND Y = 15 else
"0000000000001" when X = 36 AND Y = 15 else
"0000000000001" when X = 37 AND Y = 15 else
"0000000000001" when X = 38 AND Y = 15 else
"0000000000001" when X = 39 AND Y = 15 else
"0000000000001" when X = 40 AND Y = 15 else
"0000000000001" when X = 41 AND Y = 15 else
"0000000000001" when X = 42 AND Y = 15 else
"0111101010101" when X = 43 AND Y = 15 else
"1111111100000" when X = 44 AND Y = 15 else
"1111111100000" when X = 45 AND Y = 15 else
"1111111100000" when X = 0 AND Y = 16 else
"0101011110001" when X = 1 AND Y = 16 else
"0000000000001" when X = 2 AND Y = 16 else
"0000000000001" when X = 3 AND Y = 16 else
"0000000000001" when X = 4 AND Y = 16 else
"0000000000001" when X = 5 AND Y = 16 else
"0000000000001" when X = 6 AND Y = 16 else
"0000000000001" when X = 7 AND Y = 16 else
"0000000000001" when X = 8 AND Y = 16 else
"0000000000001" when X = 9 AND Y = 16 else
"0010000001101" when X = 10 AND Y = 16 else
"0101000110111" when X = 11 AND Y = 16 else
"0001000011111" when X = 12 AND Y = 16 else
"0000010011011" when X = 13 AND Y = 16 else
"0000100110001" when X = 14 AND Y = 16 else
"0001100010001" when X = 15 AND Y = 16 else
"0101010010011" when X = 16 AND Y = 16 else
"0111000110011" when X = 17 AND Y = 16 else
"0101010110011" when X = 18 AND Y = 16 else
"0101001110011" when X = 19 AND Y = 16 else
"1001000010001" when X = 20 AND Y = 16 else
"1111000000001" when X = 21 AND Y = 16 else
"1111000000001" when X = 22 AND Y = 16 else
"1110000000101" when X = 23 AND Y = 16 else
"1000000010001" when X = 24 AND Y = 16 else
"0101010010011" when X = 25 AND Y = 16 else
"0101010010011" when X = 26 AND Y = 16 else
"0111000010011" when X = 27 AND Y = 16 else
"0101010010011" when X = 28 AND Y = 16 else
"0001100010001" when X = 29 AND Y = 16 else
"0000100110001" when X = 30 AND Y = 16 else
"0000010011011" when X = 31 AND Y = 16 else
"0001000011111" when X = 32 AND Y = 16 else
"0101000110111" when X = 33 AND Y = 16 else
"0010000001101" when X = 34 AND Y = 16 else
"0000000000001" when X = 35 AND Y = 16 else
"0000000000001" when X = 36 AND Y = 16 else
"0000000000001" when X = 37 AND Y = 16 else
"0000000000001" when X = 38 AND Y = 16 else
"0000000000001" when X = 39 AND Y = 16 else
"0000000000001" when X = 40 AND Y = 16 else
"0000000000001" when X = 41 AND Y = 16 else
"0000000000001" when X = 42 AND Y = 16 else
"0111101010101" when X = 43 AND Y = 16 else
"1111111100000" when X = 44 AND Y = 16 else
"1111111100000" when X = 45 AND Y = 16 else
"1111111100000" when X = 0 AND Y = 17 else
"0101011110001" when X = 1 AND Y = 17 else
"0000000000001" when X = 2 AND Y = 17 else
"0000000000001" when X = 3 AND Y = 17 else
"0000000000001" when X = 4 AND Y = 17 else
"0000000000001" when X = 5 AND Y = 17 else
"0000000000001" when X = 6 AND Y = 17 else
"0000000000001" when X = 7 AND Y = 17 else
"0000000000001" when X = 8 AND Y = 17 else
"0000000000001" when X = 9 AND Y = 17 else
"0011000001001" when X = 10 AND Y = 17 else
"0101000010111" when X = 11 AND Y = 17 else
"0010001011011" when X = 12 AND Y = 17 else
"0010011010101" when X = 13 AND Y = 17 else
"0010100010011" when X = 14 AND Y = 17 else
"0011011110011" when X = 15 AND Y = 17 else
"0110001010011" when X = 16 AND Y = 17 else
"0111000010011" when X = 17 AND Y = 17 else
"0100010110011" when X = 18 AND Y = 17 else
"0110010010011" when X = 19 AND Y = 17 else
"1001001010001" when X = 20 AND Y = 17 else
"1111001000101" when X = 21 AND Y = 17 else
"1111001000011" when X = 22 AND Y = 17 else
"1110001000111" when X = 23 AND Y = 17 else
"1000001010011" when X = 24 AND Y = 17 else
"0101010110011" when X = 25 AND Y = 17 else
"0101010010011" when X = 26 AND Y = 17 else
"0111000010011" when X = 27 AND Y = 17 else
"0110001010011" when X = 28 AND Y = 17 else
"0011011110011" when X = 29 AND Y = 17 else
"0010100010011" when X = 30 AND Y = 17 else
"0010011010101" when X = 31 AND Y = 17 else
"0010001011011" when X = 32 AND Y = 17 else
"0101000010111" when X = 33 AND Y = 17 else
"0011000001001" when X = 34 AND Y = 17 else
"0000000000001" when X = 35 AND Y = 17 else
"0000000000001" when X = 36 AND Y = 17 else
"0000000000001" when X = 37 AND Y = 17 else
"0000000000001" when X = 38 AND Y = 17 else
"0000000000001" when X = 39 AND Y = 17 else
"0000000000001" when X = 40 AND Y = 17 else
"0000000000001" when X = 41 AND Y = 17 else
"0000000000001" when X = 42 AND Y = 17 else
"0111101010101" when X = 43 AND Y = 17 else
"1111111100000" when X = 44 AND Y = 17 else
"1111111100000" when X = 45 AND Y = 17 else
"1111111100000" when X = 0 AND Y = 18 else
"0110100010011" when X = 1 AND Y = 18 else
"0000000000001" when X = 2 AND Y = 18 else
"0000000000001" when X = 3 AND Y = 18 else
"0000000000001" when X = 4 AND Y = 18 else
"0000000000001" when X = 5 AND Y = 18 else
"0000000000001" when X = 6 AND Y = 18 else
"0000000000001" when X = 7 AND Y = 18 else
"0000000000001" when X = 8 AND Y = 18 else
"0000000000001" when X = 9 AND Y = 18 else
"0011000001001" when X = 10 AND Y = 18 else
"0111000010011" when X = 11 AND Y = 18 else
"0110000110101" when X = 12 AND Y = 18 else
"0110001010011" when X = 13 AND Y = 18 else
"0110001010011" when X = 14 AND Y = 18 else
"0110000110011" when X = 15 AND Y = 18 else
"0110000110011" when X = 16 AND Y = 18 else
"0111000010011" when X = 17 AND Y = 18 else
"0101010110011" when X = 18 AND Y = 18 else
"0111100110011" when X = 19 AND Y = 18 else
"1010100010011" when X = 20 AND Y = 18 else
"1010100110001" when X = 21 AND Y = 18 else
"1010100110001" when X = 22 AND Y = 18 else
"1010100010011" when X = 23 AND Y = 18 else
"1001100010011" when X = 24 AND Y = 18 else
"0110100010011" when X = 25 AND Y = 18 else
"0101010010011" when X = 26 AND Y = 18 else
"0111000010011" when X = 27 AND Y = 18 else
"0110000110011" when X = 28 AND Y = 18 else
"0110000110011" when X = 29 AND Y = 18 else
"0110001010011" when X = 30 AND Y = 18 else
"0110001010011" when X = 31 AND Y = 18 else
"0110000110101" when X = 32 AND Y = 18 else
"0111000010011" when X = 33 AND Y = 18 else
"0011000001001" when X = 34 AND Y = 18 else
"0000000000001" when X = 35 AND Y = 18 else
"0000000000001" when X = 36 AND Y = 18 else
"0000000000001" when X = 37 AND Y = 18 else
"0000000000001" when X = 38 AND Y = 18 else
"0000000000001" when X = 39 AND Y = 18 else
"0000000000001" when X = 40 AND Y = 18 else
"0000000000001" when X = 41 AND Y = 18 else
"0001000100011" when X = 42 AND Y = 18 else
"0111101010111" when X = 43 AND Y = 18 else
"1111111100000" when X = 44 AND Y = 18 else
"1111111100000" when X = 45 AND Y = 18 else
"1111111100000" when X = 0 AND Y = 19 else
"1001101111001" when X = 1 AND Y = 19 else
"0011001100111" when X = 2 AND Y = 19 else
"0000000000001" when X = 3 AND Y = 19 else
"0000000000001" when X = 4 AND Y = 19 else
"0000000000001" when X = 5 AND Y = 19 else
"0000000000001" when X = 6 AND Y = 19 else
"0000000000001" when X = 7 AND Y = 19 else
"0000000000001" when X = 8 AND Y = 19 else
"0000000000001" when X = 9 AND Y = 19 else
"0011000001001" when X = 10 AND Y = 19 else
"0110000010101" when X = 11 AND Y = 19 else
"0100000110111" when X = 12 AND Y = 19 else
"0101010010011" when X = 13 AND Y = 19 else
"0101010010011" when X = 14 AND Y = 19 else
"0101010010011" when X = 15 AND Y = 19 else
"0110000110011" when X = 16 AND Y = 19 else
"0111000010011" when X = 17 AND Y = 19 else
"0101010110011" when X = 18 AND Y = 19 else
"0111100110011" when X = 19 AND Y = 19 else
"0111100110011" when X = 20 AND Y = 19 else
"0110100110011" when X = 21 AND Y = 19 else
"0110100110011" when X = 22 AND Y = 19 else
"0110100110011" when X = 23 AND Y = 19 else
"0111100110011" when X = 24 AND Y = 19 else
"0110100110011" when X = 25 AND Y = 19 else
"0101010010011" when X = 26 AND Y = 19 else
"0111000010011" when X = 27 AND Y = 19 else
"0110000110011" when X = 28 AND Y = 19 else
"0101010010011" when X = 29 AND Y = 19 else
"0101010010011" when X = 30 AND Y = 19 else
"0101010010011" when X = 31 AND Y = 19 else
"0100000110111" when X = 32 AND Y = 19 else
"0110000010101" when X = 33 AND Y = 19 else
"0011000001001" when X = 34 AND Y = 19 else
"0000000000001" when X = 35 AND Y = 19 else
"0000000000001" when X = 36 AND Y = 19 else
"0000000000001" when X = 37 AND Y = 19 else
"0000000000001" when X = 38 AND Y = 19 else
"0000000000001" when X = 39 AND Y = 19 else
"0000000000001" when X = 40 AND Y = 19 else
"0000000000001" when X = 41 AND Y = 19 else
"0101010101011" when X = 42 AND Y = 19 else
"1110110101011" when X = 43 AND Y = 19 else
"1111111100000" when X = 44 AND Y = 19 else
"1111111100000" when X = 45 AND Y = 19 else
"1111111100000" when X = 0 AND Y = 20 else
"1001101111001" when X = 1 AND Y = 20 else
"0011001100111" when X = 2 AND Y = 20 else
"0000000000001" when X = 3 AND Y = 20 else
"0000000000001" when X = 4 AND Y = 20 else
"0000000000001" when X = 5 AND Y = 20 else
"0000000000001" when X = 6 AND Y = 20 else
"0000000000001" when X = 7 AND Y = 20 else
"0000000000001" when X = 8 AND Y = 20 else
"0000000000001" when X = 9 AND Y = 20 else
"0011000001011" when X = 10 AND Y = 20 else
"0100000111001" when X = 11 AND Y = 20 else
"0001010110111" when X = 12 AND Y = 20 else
"0000100010011" when X = 13 AND Y = 20 else
"0000100110001" when X = 14 AND Y = 20 else
"0001100010011" when X = 15 AND Y = 20 else
"0110001010011" when X = 16 AND Y = 20 else
"0110000010011" when X = 17 AND Y = 20 else
"0101010110011" when X = 18 AND Y = 20 else
"0110100110011" when X = 19 AND Y = 20 else
"0010100110011" when X = 20 AND Y = 20 else
"0000011110101" when X = 21 AND Y = 20 else
"0000010011011" when X = 22 AND Y = 20 else
"0000011110101" when X = 23 AND Y = 20 else
"0100100110011" when X = 24 AND Y = 20 else
"0110100110011" when X = 25 AND Y = 20 else
"0101010010011" when X = 26 AND Y = 20 else
"0110000010011" when X = 27 AND Y = 20 else
"0110001010011" when X = 28 AND Y = 20 else
"0001100010011" when X = 29 AND Y = 20 else
"0000100110001" when X = 30 AND Y = 20 else
"0000100010011" when X = 31 AND Y = 20 else
"0001010110111" when X = 32 AND Y = 20 else
"0100000111001" when X = 33 AND Y = 20 else
"0011000001011" when X = 34 AND Y = 20 else
"0000000000001" when X = 35 AND Y = 20 else
"0000000000001" when X = 36 AND Y = 20 else
"0000000000001" when X = 37 AND Y = 20 else
"0000000000001" when X = 38 AND Y = 20 else
"0000000000001" when X = 39 AND Y = 20 else
"0000000000001" when X = 40 AND Y = 20 else
"0000000000001" when X = 41 AND Y = 20 else
"0101010101011" when X = 42 AND Y = 20 else
"1110110101011" when X = 43 AND Y = 20 else
"1111111100000" when X = 44 AND Y = 20 else
"1111111100000" when X = 45 AND Y = 20 else
"1111111100000" when X = 0 AND Y = 21 else
"0110100010011" when X = 1 AND Y = 21 else
"0000000000001" when X = 2 AND Y = 21 else
"0000000000001" when X = 3 AND Y = 21 else
"0000000000001" when X = 4 AND Y = 21 else
"0000000000001" when X = 5 AND Y = 21 else
"0000000000001" when X = 6 AND Y = 21 else
"0000000000001" when X = 7 AND Y = 21 else
"0000000000001" when X = 8 AND Y = 21 else
"0000000000001" when X = 9 AND Y = 21 else
"0001000101111" when X = 10 AND Y = 21 else
"0001000111111" when X = 11 AND Y = 21 else
"0000011110101" when X = 12 AND Y = 21 else
"0000100110001" when X = 13 AND Y = 21 else
"0000100010011" when X = 14 AND Y = 21 else
"0000010011011" when X = 15 AND Y = 21 else
"0010000011101" when X = 16 AND Y = 21 else
"0011000011011" when X = 17 AND Y = 21 else
"0100010110011" when X = 18 AND Y = 21 else
"0110100110011" when X = 19 AND Y = 21 else
"0010100110011" when X = 20 AND Y = 21 else
"0000011010111" when X = 21 AND Y = 21 else
"0001001011111" when X = 22 AND Y = 21 else
"0000011110101" when X = 23 AND Y = 21 else
"0100100110011" when X = 24 AND Y = 21 else
"0110100110011" when X = 25 AND Y = 21 else
"0101010010011" when X = 26 AND Y = 21 else
"0011000011011" when X = 27 AND Y = 21 else
"0010000011101" when X = 28 AND Y = 21 else
"0000010011011" when X = 29 AND Y = 21 else
"0000100010011" when X = 30 AND Y = 21 else
"0000100110001" when X = 31 AND Y = 21 else
"0000011110101" when X = 32 AND Y = 21 else
"0001000111111" when X = 33 AND Y = 21 else
"0001000101111" when X = 34 AND Y = 21 else
"0000000000001" when X = 35 AND Y = 21 else
"0000000000001" when X = 36 AND Y = 21 else
"0000000000001" when X = 37 AND Y = 21 else
"0000000000001" when X = 38 AND Y = 21 else
"0000000000001" when X = 39 AND Y = 21 else
"0000000000001" when X = 40 AND Y = 21 else
"0000000000001" when X = 41 AND Y = 21 else
"0001000100011" when X = 42 AND Y = 21 else
"0111101010111" when X = 43 AND Y = 21 else
"1111111100000" when X = 44 AND Y = 21 else
"1111111100000" when X = 45 AND Y = 21 else
"1111111100000" when X = 0 AND Y = 22 else
"0101011110001" when X = 1 AND Y = 22 else
"0000000000001" when X = 2 AND Y = 22 else
"0000000000001" when X = 3 AND Y = 22 else
"0000000000001" when X = 4 AND Y = 22 else
"0000000000001" when X = 5 AND Y = 22 else
"0000000000001" when X = 6 AND Y = 22 else
"0000000000001" when X = 7 AND Y = 22 else
"0000000000001" when X = 8 AND Y = 22 else
"0000000000001" when X = 9 AND Y = 22 else
"0100010101111" when X = 10 AND Y = 22 else
"0100011111111" when X = 11 AND Y = 22 else
"0000001111101" when X = 12 AND Y = 22 else
"0000011110101" when X = 13 AND Y = 22 else
"0000010111001" when X = 14 AND Y = 22 else
"0001000011111" when X = 15 AND Y = 22 else
"0001000011111" when X = 16 AND Y = 22 else
"0001000011111" when X = 17 AND Y = 22 else
"0001010110111" when X = 18 AND Y = 22 else
"0111100110011" when X = 19 AND Y = 22 else
"0010100110011" when X = 20 AND Y = 22 else
"0000100010011" when X = 21 AND Y = 22 else
"0000100010011" when X = 22 AND Y = 22 else
"0000100010011" when X = 23 AND Y = 22 else
"0100100110011" when X = 24 AND Y = 22 else
"0110100110011" when X = 25 AND Y = 22 else
"0001010011001" when X = 26 AND Y = 22 else
"0001000011111" when X = 27 AND Y = 22 else
"0001000011111" when X = 28 AND Y = 22 else
"0001000011111" when X = 29 AND Y = 22 else
"0000010111001" when X = 30 AND Y = 22 else
"0000011110101" when X = 31 AND Y = 22 else
"0000001111101" when X = 32 AND Y = 22 else
"0100011111111" when X = 33 AND Y = 22 else
"0100011001111" when X = 34 AND Y = 22 else
"0000000000001" when X = 35 AND Y = 22 else
"0000000000001" when X = 36 AND Y = 22 else
"0000000000001" when X = 37 AND Y = 22 else
"0000000000001" when X = 38 AND Y = 22 else
"0000000000001" when X = 39 AND Y = 22 else
"0000000000001" when X = 40 AND Y = 22 else
"0000000000001" when X = 41 AND Y = 22 else
"0000000000001" when X = 42 AND Y = 22 else
"0111101010101" when X = 43 AND Y = 22 else
"1111111100000" when X = 44 AND Y = 22 else
"1111111100000" when X = 45 AND Y = 22 else
"1111111100000" when X = 0 AND Y = 23 else
"0101011110001" when X = 1 AND Y = 23 else
"0000000000001" when X = 2 AND Y = 23 else
"0000000000001" when X = 3 AND Y = 23 else
"0000000000001" when X = 4 AND Y = 23 else
"0000000000001" when X = 5 AND Y = 23 else
"0000000000001" when X = 6 AND Y = 23 else
"0000000000001" when X = 7 AND Y = 23 else
"0000000000001" when X = 8 AND Y = 23 else
"0000000000001" when X = 9 AND Y = 23 else
"0100011001111" when X = 10 AND Y = 23 else
"1111111100000" when X = 11 AND Y = 23 else
"0100011011111" when X = 12 AND Y = 23 else
"0000001111101" when X = 13 AND Y = 23 else
"0000001111101" when X = 14 AND Y = 23 else
"0001000011111" when X = 15 AND Y = 23 else
"0001000011111" when X = 16 AND Y = 23 else
"0001000011111" when X = 17 AND Y = 23 else
"0000010111001" when X = 18 AND Y = 23 else
"0111100110011" when X = 19 AND Y = 23 else
"0110100110011" when X = 20 AND Y = 23 else
"0101100110011" when X = 21 AND Y = 23 else
"0101100110011" when X = 22 AND Y = 23 else
"0101100110011" when X = 23 AND Y = 23 else
"0110100110011" when X = 24 AND Y = 23 else
"0110100110011" when X = 25 AND Y = 23 else
"0000010011011" when X = 26 AND Y = 23 else
"0001000011111" when X = 27 AND Y = 23 else
"0001000011111" when X = 28 AND Y = 23 else
"0001000011111" when X = 29 AND Y = 23 else
"0000001111101" when X = 30 AND Y = 23 else
"0000001111101" when X = 31 AND Y = 23 else
"0011011011111" when X = 32 AND Y = 23 else
"1111111100000" when X = 33 AND Y = 23 else
"0100011001111" when X = 34 AND Y = 23 else
"0000000000001" when X = 35 AND Y = 23 else
"0000000000001" when X = 36 AND Y = 23 else
"0000000000001" when X = 37 AND Y = 23 else
"0000000000001" when X = 38 AND Y = 23 else
"0000000000001" when X = 39 AND Y = 23 else
"0000000000001" when X = 40 AND Y = 23 else
"0000000000001" when X = 41 AND Y = 23 else
"0000000000001" when X = 42 AND Y = 23 else
"0111101010101" when X = 43 AND Y = 23 else
"1111111100000" when X = 44 AND Y = 23 else
"1111111100000" when X = 45 AND Y = 23 else
"1111111100000" when X = 0 AND Y = 24 else
"0101100010001" when X = 1 AND Y = 24 else
"0000000000001" when X = 2 AND Y = 24 else
"0000000000001" when X = 3 AND Y = 24 else
"0000000000001" when X = 4 AND Y = 24 else
"0000000000001" when X = 5 AND Y = 24 else
"0000000000001" when X = 6 AND Y = 24 else
"0000000000001" when X = 7 AND Y = 24 else
"0000000000001" when X = 8 AND Y = 24 else
"0000000000001" when X = 9 AND Y = 24 else
"0100011001111" when X = 10 AND Y = 24 else
"1111111100000" when X = 11 AND Y = 24 else
"1111111100000" when X = 12 AND Y = 24 else
"0101100111111" when X = 13 AND Y = 24 else
"0101100011111" when X = 14 AND Y = 24 else
"0010001111111" when X = 15 AND Y = 24 else
"0001000011111" when X = 16 AND Y = 24 else
"0010010011111" when X = 17 AND Y = 24 else
"0110101011011" when X = 18 AND Y = 24 else
"1000110011001" when X = 19 AND Y = 24 else
"1001110011001" when X = 20 AND Y = 24 else
"1001110011001" when X = 21 AND Y = 24 else
"1001110011001" when X = 22 AND Y = 24 else
"1001110011001" when X = 23 AND Y = 24 else
"1001110011001" when X = 24 AND Y = 24 else
"1000101111001" when X = 25 AND Y = 24 else
"0101100111101" when X = 26 AND Y = 24 else
"0010010011111" when X = 27 AND Y = 24 else
"0001000011111" when X = 28 AND Y = 24 else
"0010001111111" when X = 29 AND Y = 24 else
"0101100011111" when X = 30 AND Y = 24 else
"0101100111111" when X = 31 AND Y = 24 else
"1111111100000" when X = 32 AND Y = 24 else
"1111111100000" when X = 33 AND Y = 24 else
"0100011101111" when X = 34 AND Y = 24 else
"0000000000001" when X = 35 AND Y = 24 else
"0000000000001" when X = 36 AND Y = 24 else
"0000000000001" when X = 37 AND Y = 24 else
"0000000000001" when X = 38 AND Y = 24 else
"0000000000001" when X = 39 AND Y = 24 else
"0000000000001" when X = 40 AND Y = 24 else
"0000000000001" when X = 41 AND Y = 24 else
"0000000000001" when X = 42 AND Y = 24 else
"0111101010101" when X = 43 AND Y = 24 else
"1111111100000" when X = 44 AND Y = 24 else
"1111111100000" when X = 45 AND Y = 24 else
"1111111100000" when X = 0 AND Y = 25 else
"1000110011011" when X = 1 AND Y = 25 else
"0011010101011" when X = 2 AND Y = 25 else
"0001000100011" when X = 3 AND Y = 25 else
"0001000100011" when X = 4 AND Y = 25 else
"0001000100011" when X = 5 AND Y = 25 else
"0001000100011" when X = 6 AND Y = 25 else
"0001000100011" when X = 7 AND Y = 25 else
"0001000100011" when X = 8 AND Y = 25 else
"0011010001001" when X = 9 AND Y = 25 else
"1000101111001" when X = 10 AND Y = 25 else
"1111111100000" when X = 11 AND Y = 25 else
"1111111100000" when X = 12 AND Y = 25 else
"1111111100000" when X = 13 AND Y = 25 else
"1111111100000" when X = 14 AND Y = 25 else
"0111101111101" when X = 15 AND Y = 25 else
"0110101011111" when X = 16 AND Y = 25 else
"1000101111101" when X = 17 AND Y = 25 else
"1111111100000" when X = 18 AND Y = 25 else
"1111111100000" when X = 19 AND Y = 25 else
"1111111100000" when X = 20 AND Y = 25 else
"1111111100000" when X = 21 AND Y = 25 else
"1111111100000" when X = 22 AND Y = 25 else
"1111111100000" when X = 23 AND Y = 25 else
"1111111100000" when X = 24 AND Y = 25 else
"1111111100000" when X = 25 AND Y = 25 else
"1111111100000" when X = 26 AND Y = 25 else
"1000101111101" when X = 27 AND Y = 25 else
"0110101011111" when X = 28 AND Y = 25 else
"0111101111101" when X = 29 AND Y = 25 else
"1111111100000" when X = 30 AND Y = 25 else
"1111111100000" when X = 31 AND Y = 25 else
"1111111100000" when X = 32 AND Y = 25 else
"1111111100000" when X = 33 AND Y = 25 else
"1000101111001" when X = 34 AND Y = 25 else
"0011010001001" when X = 35 AND Y = 25 else
"0001000100011" when X = 36 AND Y = 25 else
"0001000100011" when X = 37 AND Y = 25 else
"0001000100011" when X = 38 AND Y = 25 else
"0001000100011" when X = 39 AND Y = 25 else
"0001000100011" when X = 40 AND Y = 25 else
"0001000100011" when X = 41 AND Y = 25 else
"0100011001111" when X = 42 AND Y = 25 else
"1111111100000" when X = 43 AND Y = 25 else
"1111111100000" when X = 44 AND Y = 25 else
"1111111100000" when X = 45 AND Y = 25 else
"1111111100000" when X = 0 AND Y = 26 else
"1111111100000" when X = 1 AND Y = 26 else
"1111111100000" when X = 2 AND Y = 26 else
"1000101111001" when X = 3 AND Y = 26 else
"1000101111001" when X = 4 AND Y = 26 else
"1000101111001" when X = 5 AND Y = 26 else
"1000101111001" when X = 6 AND Y = 26 else
"1000101111001" when X = 7 AND Y = 26 else
"1000101111001" when X = 8 AND Y = 26 else
"1110110101001" when X = 9 AND Y = 26 else
"1111111100000" when X = 10 AND Y = 26 else
"1111111100000" when X = 11 AND Y = 26 else
"1111111100000" when X = 12 AND Y = 26 else
"1111111100000" when X = 13 AND Y = 26 else
"1111111100000" when X = 14 AND Y = 26 else
"1111111100000" when X = 15 AND Y = 26 else
"1111111100000" when X = 16 AND Y = 26 else
"1111111100000" when X = 17 AND Y = 26 else
"1111111100000" when X = 18 AND Y = 26 else
"1111111100000" when X = 19 AND Y = 26 else
"1111111100000" when X = 20 AND Y = 26 else
"1111111100000" when X = 21 AND Y = 26 else
"1111111100000" when X = 22 AND Y = 26 else
"1111111100000" when X = 23 AND Y = 26 else
"1111111100000" when X = 24 AND Y = 26 else
"1111111100000" when X = 25 AND Y = 26 else
"1111111100000" when X = 26 AND Y = 26 else
"1111111100000" when X = 27 AND Y = 26 else
"1111111100000" when X = 28 AND Y = 26 else
"1111111100000" when X = 29 AND Y = 26 else
"1111111100000" when X = 30 AND Y = 26 else
"1111111100000" when X = 31 AND Y = 26 else
"1111111100000" when X = 32 AND Y = 26 else
"1111111100000" when X = 33 AND Y = 26 else
"1111111100000" when X = 34 AND Y = 26 else
"1110110101001" when X = 35 AND Y = 26 else
"1000101111001" when X = 36 AND Y = 26 else
"1000101111001" when X = 37 AND Y = 26 else
"1000101111001" when X = 38 AND Y = 26 else
"1000101111001" when X = 39 AND Y = 26 else
"1000101111001" when X = 40 AND Y = 26 else
"1000101111001" when X = 41 AND Y = 26 else
"1111111100000" when X = 42 AND Y = 26 else
"1111111100000" when X = 43 AND Y = 26 else
"1111111100000" when X = 44 AND Y = 26 else
"1111111100000" when X = 45 AND Y = 26 else
"1111111100000" when X = 0 AND Y = 27 else
"1111111100000" when X = 1 AND Y = 27 else
"1111111100000" when X = 2 AND Y = 27 else
"1111111100000" when X = 3 AND Y = 27 else
"1111111100000" when X = 4 AND Y = 27 else
"1111111100000" when X = 5 AND Y = 27 else
"1111111100000" when X = 6 AND Y = 27 else
"1111111100000" when X = 7 AND Y = 27 else
"1111111100000" when X = 8 AND Y = 27 else
"1111111100000" when X = 9 AND Y = 27 else
"1111111100000" when X = 10 AND Y = 27 else
"1111111100000" when X = 11 AND Y = 27 else
"1111111100000" when X = 12 AND Y = 27 else
"1111111100000" when X = 13 AND Y = 27 else
"1111111100000" when X = 14 AND Y = 27 else
"1111111100000" when X = 15 AND Y = 27 else
"1111111100000" when X = 16 AND Y = 27 else
"1111111100000" when X = 17 AND Y = 27 else
"1111111100000" when X = 18 AND Y = 27 else
"1111111100000" when X = 19 AND Y = 27 else
"1111111100000" when X = 20 AND Y = 27 else
"1111111100000" when X = 21 AND Y = 27 else
"1111111100000" when X = 22 AND Y = 27 else
"1111111100000" when X = 23 AND Y = 27 else
"1111111100000" when X = 24 AND Y = 27 else
"1111111100000" when X = 25 AND Y = 27 else
"1111111100000" when X = 26 AND Y = 27 else
"1111111100000" when X = 27 AND Y = 27 else
"1111111100000" when X = 28 AND Y = 27 else
"1111111100000" when X = 29 AND Y = 27 else
"1111111100000" when X = 30 AND Y = 27 else
"1111111100000" when X = 31 AND Y = 27 else
"1111111100000" when X = 32 AND Y = 27 else
"1111111100000" when X = 33 AND Y = 27 else
"1111111100000" when X = 34 AND Y = 27 else
"1111111100000" when X = 35 AND Y = 27 else
"1111111100000" when X = 36 AND Y = 27 else
"1111111100000" when X = 37 AND Y = 27 else
"1111111100000" when X = 38 AND Y = 27 else
"1111111100000" when X = 39 AND Y = 27 else
"1111111100000" when X = 40 AND Y = 27 else
"1111111100000" when X = 41 AND Y = 27 else
"1111111100000" when X = 42 AND Y = 27 else
"1111111100000" when X = 43 AND Y = 27 else
"1111111100000" when X = 44 AND Y = 27 else
"1111111100000" when X = 45 AND Y = 27 else
"1111111100000" when X = 0 AND Y = 28 else
"1111111100000" when X = 1 AND Y = 28 else
"1111111100000" when X = 2 AND Y = 28 else
"1111111100000" when X = 3 AND Y = 28 else
"1111111100000" when X = 4 AND Y = 28 else
"1111111100000" when X = 5 AND Y = 28 else
"1111111100000" when X = 6 AND Y = 28 else
"1111111100000" when X = 7 AND Y = 28 else
"1111111100000" when X = 8 AND Y = 28 else
"1111111100000" when X = 9 AND Y = 28 else
"1111111100000" when X = 10 AND Y = 28 else
"1111111100000" when X = 11 AND Y = 28 else
"1111111100000" when X = 12 AND Y = 28 else
"1111111100000" when X = 13 AND Y = 28 else
"1111111100000" when X = 14 AND Y = 28 else
"1111111100000" when X = 15 AND Y = 28 else
"1111111100000" when X = 16 AND Y = 28 else
"1111111100000" when X = 17 AND Y = 28 else
"1111111100000" when X = 18 AND Y = 28 else
"1111111100000" when X = 19 AND Y = 28 else
"1111111100000" when X = 20 AND Y = 28 else
"1111111100000" when X = 21 AND Y = 28 else
"1111111100000" when X = 22 AND Y = 28 else
"1111111100000" when X = 23 AND Y = 28 else
"1111111100000" when X = 24 AND Y = 28 else
"1111111100000" when X = 25 AND Y = 28 else
"1111111100000" when X = 26 AND Y = 28 else
"1111111100000" when X = 27 AND Y = 28 else
"1111111100000" when X = 28 AND Y = 28 else
"1111111100000" when X = 29 AND Y = 28 else
"1111111100000" when X = 30 AND Y = 28 else
"1111111100000" when X = 31 AND Y = 28 else
"1111111100000" when X = 32 AND Y = 28 else
"1111111100000" when X = 33 AND Y = 28 else
"1111111100000" when X = 34 AND Y = 28 else
"1111111100000" when X = 35 AND Y = 28 else
"1111111100000" when X = 36 AND Y = 28 else
"1111111100000" when X = 37 AND Y = 28 else
"1111111100000" when X = 38 AND Y = 28 else
"1111111100000" when X = 39 AND Y = 28 else
"1111111100000" when X = 40 AND Y = 28 else
"1111111100000" when X = 41 AND Y = 28 else
"1111111100000" when X = 42 AND Y = 28 else
"1111111100000" when X = 43 AND Y = 28 else
"1111111100000" when X = 44 AND Y = 28 else
"1111111100000" when X = 45 AND Y = 28 else
"1111111100000" when X = 0 AND Y = 29 else
"1111111100000" when X = 1 AND Y = 29 else
"1111111100000" when X = 2 AND Y = 29 else
"1111111100000" when X = 3 AND Y = 29 else
"1111111100000" when X = 4 AND Y = 29 else
"1111111100000" when X = 5 AND Y = 29 else
"1111111100000" when X = 6 AND Y = 29 else
"1111111100000" when X = 7 AND Y = 29 else
"1111111100000" when X = 8 AND Y = 29 else
"1111111100000" when X = 9 AND Y = 29 else
"1111111100000" when X = 10 AND Y = 29 else
"1111111100000" when X = 11 AND Y = 29 else
"1111111100000" when X = 12 AND Y = 29 else
"1111111100000" when X = 13 AND Y = 29 else
"1111111100000" when X = 14 AND Y = 29 else
"1111111100000" when X = 15 AND Y = 29 else
"1111111100000" when X = 16 AND Y = 29 else
"1111111100000" when X = 17 AND Y = 29 else
"1111111100000" when X = 18 AND Y = 29 else
"1111111100000" when X = 19 AND Y = 29 else
"1111111100000" when X = 20 AND Y = 29 else
"1111111100000" when X = 21 AND Y = 29 else
"1111111100000" when X = 22 AND Y = 29 else
"1111111100000" when X = 23 AND Y = 29 else
"1111111100000" when X = 24 AND Y = 29 else
"1111111100000" when X = 25 AND Y = 29 else
"1111111100000" when X = 26 AND Y = 29 else
"1111111100000" when X = 27 AND Y = 29 else
"1111111100000" when X = 28 AND Y = 29 else
"1111111100000" when X = 29 AND Y = 29 else
"1111111100000" when X = 30 AND Y = 29 else
"1111111100000" when X = 31 AND Y = 29 else
"1111111100000" when X = 32 AND Y = 29 else
"1111111100000" when X = 33 AND Y = 29 else
"1111111100000" when X = 34 AND Y = 29 else
"1111111100000" when X = 35 AND Y = 29 else
"1111111100000" when X = 36 AND Y = 29 else
"1111111100000" when X = 37 AND Y = 29 else
"1111111100000" when X = 38 AND Y = 29 else
"1111111100000" when X = 39 AND Y = 29 else
"1111111100000" when X = 40 AND Y = 29 else
"1111111100000" when X = 41 AND Y = 29 else
"1111111100000" when X = 42 AND Y = 29 else
"1111111100000" when X = 43 AND Y = 29 else
"1111111100000" when X = 44 AND Y = 29 else
"1111111100000" when X = 45 AND Y = 29 else
"0000000000000"; -- should never get here
end rtl;
