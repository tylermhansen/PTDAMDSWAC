-- Tyler Hansen
-- CS232 Final Project
-- genSpriteROM.py
-- generates a ROM file in VHDL from a .ppm image

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity player_sprite_straight_updated is
port(
X	: in INTEGER RANGE 0 TO 1688;
Y	: in INTEGER RANGE 0 TO 1688;
data : out std_logic_vector (11 downto 0)
);

end entity;

architecture rtl of player_sprite_straight_updated is
begin
data <=
"111111110000" when X = 0 AND Y = 0 else
"111111110000" when X = 1 AND Y = 0 else
"111111110000" when X = 2 AND Y = 0 else
"111111110000" when X = 3 AND Y = 0 else
"111111110000" when X = 4 AND Y = 0 else
"111111110000" when X = 5 AND Y = 0 else
"111111110000" when X = 6 AND Y = 0 else
"111111110000" when X = 7 AND Y = 0 else
"111111110000" when X = 8 AND Y = 0 else
"111111110000" when X = 9 AND Y = 0 else
"111111110000" when X = 10 AND Y = 0 else
"111111110000" when X = 11 AND Y = 0 else
"111111110000" when X = 12 AND Y = 0 else
"111111110000" when X = 13 AND Y = 0 else
"111111110000" when X = 14 AND Y = 0 else
"111111110000" when X = 15 AND Y = 0 else
"111111110000" when X = 16 AND Y = 0 else
"111111110000" when X = 17 AND Y = 0 else
"111111110000" when X = 18 AND Y = 0 else
"111111110000" when X = 19 AND Y = 0 else
"111111110000" when X = 20 AND Y = 0 else
"111111110000" when X = 21 AND Y = 0 else
"111111110000" when X = 22 AND Y = 0 else
"111111110000" when X = 23 AND Y = 0 else
"111111110000" when X = 24 AND Y = 0 else
"111111110000" when X = 25 AND Y = 0 else
"111111110000" when X = 26 AND Y = 0 else
"111111110000" when X = 27 AND Y = 0 else
"111111110000" when X = 28 AND Y = 0 else
"111111110000" when X = 29 AND Y = 0 else
"111111110000" when X = 30 AND Y = 0 else
"111111110000" when X = 31 AND Y = 0 else
"111111110000" when X = 32 AND Y = 0 else
"111111110000" when X = 33 AND Y = 0 else
"111111110000" when X = 34 AND Y = 0 else
"111111110000" when X = 35 AND Y = 0 else
"111111110000" when X = 36 AND Y = 0 else
"111111110000" when X = 37 AND Y = 0 else
"111111110000" when X = 38 AND Y = 0 else
"111111110000" when X = 39 AND Y = 0 else
"111111110000" when X = 40 AND Y = 0 else
"111111110000" when X = 41 AND Y = 0 else
"111111110000" when X = 42 AND Y = 0 else
"111111110000" when X = 43 AND Y = 0 else
"111111110000" when X = 44 AND Y = 0 else
"111111110000" when X = 45 AND Y = 0 else
"111111110000" when X = 0 AND Y = 1 else
"111111110000" when X = 1 AND Y = 1 else
"111111110000" when X = 2 AND Y = 1 else
"111111110000" when X = 3 AND Y = 1 else
"111111110000" when X = 4 AND Y = 1 else
"111111110000" when X = 5 AND Y = 1 else
"111111110000" when X = 6 AND Y = 1 else
"111111110000" when X = 7 AND Y = 1 else
"111111110000" when X = 8 AND Y = 1 else
"111111110000" when X = 9 AND Y = 1 else
"111111110000" when X = 10 AND Y = 1 else
"111111110000" when X = 11 AND Y = 1 else
"111111110000" when X = 12 AND Y = 1 else
"111111110000" when X = 13 AND Y = 1 else
"111111110000" when X = 14 AND Y = 1 else
"111111110000" when X = 15 AND Y = 1 else
"111111110000" when X = 16 AND Y = 1 else
"111111110000" when X = 17 AND Y = 1 else
"111111110000" when X = 18 AND Y = 1 else
"111111110000" when X = 19 AND Y = 1 else
"111111110000" when X = 20 AND Y = 1 else
"111111110000" when X = 21 AND Y = 1 else
"111111110000" when X = 22 AND Y = 1 else
"111111110000" when X = 23 AND Y = 1 else
"111111110000" when X = 24 AND Y = 1 else
"111111110000" when X = 25 AND Y = 1 else
"111111110000" when X = 26 AND Y = 1 else
"111111110000" when X = 27 AND Y = 1 else
"111111110000" when X = 28 AND Y = 1 else
"111111110000" when X = 29 AND Y = 1 else
"111111110000" when X = 30 AND Y = 1 else
"111111110000" when X = 31 AND Y = 1 else
"111111110000" when X = 32 AND Y = 1 else
"111111110000" when X = 33 AND Y = 1 else
"111111110000" when X = 34 AND Y = 1 else
"111111110000" when X = 35 AND Y = 1 else
"111111110000" when X = 36 AND Y = 1 else
"111111110000" when X = 37 AND Y = 1 else
"111111110000" when X = 38 AND Y = 1 else
"111111110000" when X = 39 AND Y = 1 else
"111111110000" when X = 40 AND Y = 1 else
"111111110000" when X = 41 AND Y = 1 else
"111111110000" when X = 42 AND Y = 1 else
"111111110000" when X = 43 AND Y = 1 else
"111111110000" when X = 44 AND Y = 1 else
"111111110000" when X = 45 AND Y = 1 else
"111111110000" when X = 0 AND Y = 2 else
"111111110000" when X = 1 AND Y = 2 else
"111111110000" when X = 2 AND Y = 2 else
"111111110000" when X = 3 AND Y = 2 else
"111111110000" when X = 4 AND Y = 2 else
"111111110000" when X = 5 AND Y = 2 else
"111111110000" when X = 6 AND Y = 2 else
"111111110000" when X = 7 AND Y = 2 else
"111111110000" when X = 8 AND Y = 2 else
"111111110000" when X = 9 AND Y = 2 else
"111111110000" when X = 10 AND Y = 2 else
"111111110000" when X = 11 AND Y = 2 else
"111111110000" when X = 12 AND Y = 2 else
"111111110000" when X = 13 AND Y = 2 else
"111111110000" when X = 14 AND Y = 2 else
"111111110000" when X = 15 AND Y = 2 else
"111111110000" when X = 16 AND Y = 2 else
"111111110000" when X = 17 AND Y = 2 else
"111111110000" when X = 18 AND Y = 2 else
"111111110000" when X = 19 AND Y = 2 else
"111111110000" when X = 20 AND Y = 2 else
"111111110000" when X = 21 AND Y = 2 else
"111111110000" when X = 22 AND Y = 2 else
"111111110000" when X = 23 AND Y = 2 else
"111111110000" when X = 24 AND Y = 2 else
"111111110000" when X = 25 AND Y = 2 else
"111111110000" when X = 26 AND Y = 2 else
"111111110000" when X = 27 AND Y = 2 else
"111111110000" when X = 28 AND Y = 2 else
"111111110000" when X = 29 AND Y = 2 else
"111111110000" when X = 30 AND Y = 2 else
"111111110000" when X = 31 AND Y = 2 else
"111111110000" when X = 32 AND Y = 2 else
"111111110000" when X = 33 AND Y = 2 else
"111111110000" when X = 34 AND Y = 2 else
"111111110000" when X = 35 AND Y = 2 else
"111111110000" when X = 36 AND Y = 2 else
"111111110000" when X = 37 AND Y = 2 else
"111111110000" when X = 38 AND Y = 2 else
"111111110000" when X = 39 AND Y = 2 else
"111111110000" when X = 40 AND Y = 2 else
"111111110000" when X = 41 AND Y = 2 else
"111111110000" when X = 42 AND Y = 2 else
"111111110000" when X = 43 AND Y = 2 else
"111111110000" when X = 44 AND Y = 2 else
"111111110000" when X = 45 AND Y = 2 else
"111111110000" when X = 0 AND Y = 3 else
"111111110000" when X = 1 AND Y = 3 else
"111111110000" when X = 2 AND Y = 3 else
"111111110000" when X = 3 AND Y = 3 else
"111111110000" when X = 4 AND Y = 3 else
"111111110000" when X = 5 AND Y = 3 else
"111111110000" when X = 6 AND Y = 3 else
"111111110000" when X = 7 AND Y = 3 else
"111111110000" when X = 8 AND Y = 3 else
"111111110000" when X = 9 AND Y = 3 else
"111111110000" when X = 10 AND Y = 3 else
"111111110000" when X = 11 AND Y = 3 else
"111111110000" when X = 12 AND Y = 3 else
"111111110000" when X = 13 AND Y = 3 else
"111111110000" when X = 14 AND Y = 3 else
"111111110000" when X = 15 AND Y = 3 else
"111111110000" when X = 16 AND Y = 3 else
"111111110000" when X = 17 AND Y = 3 else
"111111110000" when X = 18 AND Y = 3 else
"111111110000" when X = 19 AND Y = 3 else
"011110111110" when X = 20 AND Y = 3 else
"010001101111" when X = 21 AND Y = 3 else
"010001101111" when X = 22 AND Y = 3 else
"010001111111" when X = 23 AND Y = 3 else
"111111110000" when X = 24 AND Y = 3 else
"111111110000" when X = 25 AND Y = 3 else
"111111110000" when X = 26 AND Y = 3 else
"111111110000" when X = 27 AND Y = 3 else
"111111110000" when X = 28 AND Y = 3 else
"111111110000" when X = 29 AND Y = 3 else
"111111110000" when X = 30 AND Y = 3 else
"111111110000" when X = 31 AND Y = 3 else
"111111110000" when X = 32 AND Y = 3 else
"111111110000" when X = 33 AND Y = 3 else
"111111110000" when X = 34 AND Y = 3 else
"111111110000" when X = 35 AND Y = 3 else
"111111110000" when X = 36 AND Y = 3 else
"111111110000" when X = 37 AND Y = 3 else
"111111110000" when X = 38 AND Y = 3 else
"111111110000" when X = 39 AND Y = 3 else
"111111110000" when X = 40 AND Y = 3 else
"111111110000" when X = 41 AND Y = 3 else
"111111110000" when X = 42 AND Y = 3 else
"111111110000" when X = 43 AND Y = 3 else
"111111110000" when X = 44 AND Y = 3 else
"111111110000" when X = 45 AND Y = 3 else
"111111110000" when X = 0 AND Y = 4 else
"111111110000" when X = 1 AND Y = 4 else
"111111110000" when X = 2 AND Y = 4 else
"111111110000" when X = 3 AND Y = 4 else
"111111110000" when X = 4 AND Y = 4 else
"111111110000" when X = 5 AND Y = 4 else
"111111110000" when X = 6 AND Y = 4 else
"111111110000" when X = 7 AND Y = 4 else
"111111110000" when X = 8 AND Y = 4 else
"111111110000" when X = 9 AND Y = 4 else
"111111110000" when X = 10 AND Y = 4 else
"111111110000" when X = 11 AND Y = 4 else
"111111110000" when X = 12 AND Y = 4 else
"111111110000" when X = 13 AND Y = 4 else
"111111110000" when X = 14 AND Y = 4 else
"111111110000" when X = 15 AND Y = 4 else
"111111110000" when X = 16 AND Y = 4 else
"111111110000" when X = 17 AND Y = 4 else
"111111110000" when X = 18 AND Y = 4 else
"100010111110" when X = 19 AND Y = 4 else
"001001011111" when X = 20 AND Y = 4 else
"001001011111" when X = 21 AND Y = 4 else
"010110101111" when X = 22 AND Y = 4 else
"000101001111" when X = 23 AND Y = 4 else
"001101101111" when X = 24 AND Y = 4 else
"111111110000" when X = 25 AND Y = 4 else
"111111110000" when X = 26 AND Y = 4 else
"111111110000" when X = 27 AND Y = 4 else
"111111110000" when X = 28 AND Y = 4 else
"111111110000" when X = 29 AND Y = 4 else
"111111110000" when X = 30 AND Y = 4 else
"111111110000" when X = 31 AND Y = 4 else
"111111110000" when X = 32 AND Y = 4 else
"111111110000" when X = 33 AND Y = 4 else
"111111110000" when X = 34 AND Y = 4 else
"111111110000" when X = 35 AND Y = 4 else
"111111110000" when X = 36 AND Y = 4 else
"111111110000" when X = 37 AND Y = 4 else
"111111110000" when X = 38 AND Y = 4 else
"111111110000" when X = 39 AND Y = 4 else
"111111110000" when X = 40 AND Y = 4 else
"111111110000" when X = 41 AND Y = 4 else
"111111110000" when X = 42 AND Y = 4 else
"111111110000" when X = 43 AND Y = 4 else
"111111110000" when X = 44 AND Y = 4 else
"111111110000" when X = 45 AND Y = 4 else
"111111110000" when X = 0 AND Y = 5 else
"111111110000" when X = 1 AND Y = 5 else
"111111110000" when X = 2 AND Y = 5 else
"111111110000" when X = 3 AND Y = 5 else
"111111110000" when X = 4 AND Y = 5 else
"111111110000" when X = 5 AND Y = 5 else
"111111110000" when X = 6 AND Y = 5 else
"011110101011" when X = 7 AND Y = 5 else
"011110101010" when X = 8 AND Y = 5 else
"011110101011" when X = 9 AND Y = 5 else
"100011001100" when X = 10 AND Y = 5 else
"111111110000" when X = 11 AND Y = 5 else
"111111110000" when X = 12 AND Y = 5 else
"111111110000" when X = 13 AND Y = 5 else
"111111110000" when X = 14 AND Y = 5 else
"111111110000" when X = 15 AND Y = 5 else
"101111001100" when X = 16 AND Y = 5 else
"101110111011" when X = 17 AND Y = 5 else
"100111001101" when X = 18 AND Y = 5 else
"001001011111" when X = 19 AND Y = 5 else
"000100111110" when X = 20 AND Y = 5 else
"011011001011" when X = 21 AND Y = 5 else
"011111011010" when X = 22 AND Y = 5 else
"010110111011" when X = 23 AND Y = 5 else
"000100101111" when X = 24 AND Y = 5 else
"001101111111" when X = 25 AND Y = 5 else
"101011001100" when X = 26 AND Y = 5 else
"101110111011" when X = 27 AND Y = 5 else
"101111001100" when X = 28 AND Y = 5 else
"111111110000" when X = 29 AND Y = 5 else
"111111110000" when X = 30 AND Y = 5 else
"111111110000" when X = 31 AND Y = 5 else
"111111110000" when X = 32 AND Y = 5 else
"111111110000" when X = 33 AND Y = 5 else
"100011001100" when X = 34 AND Y = 5 else
"011110101010" when X = 35 AND Y = 5 else
"011110101010" when X = 36 AND Y = 5 else
"011110111100" when X = 37 AND Y = 5 else
"111111110000" when X = 38 AND Y = 5 else
"111111110000" when X = 39 AND Y = 5 else
"111111110000" when X = 40 AND Y = 5 else
"111111110000" when X = 41 AND Y = 5 else
"111111110000" when X = 42 AND Y = 5 else
"111111110000" when X = 43 AND Y = 5 else
"111111110000" when X = 44 AND Y = 5 else
"111111110000" when X = 45 AND Y = 5 else
"111111110000" when X = 0 AND Y = 6 else
"111111110000" when X = 1 AND Y = 6 else
"111111110000" when X = 2 AND Y = 6 else
"111111110000" when X = 3 AND Y = 6 else
"111111110000" when X = 4 AND Y = 6 else
"111111110000" when X = 5 AND Y = 6 else
"011110011010" when X = 6 AND Y = 6 else
"010001010101" when X = 7 AND Y = 6 else
"001100110011" when X = 8 AND Y = 6 else
"000000000000" when X = 9 AND Y = 6 else
"001001000100" when X = 10 AND Y = 6 else
"100010111100" when X = 11 AND Y = 6 else
"111111110000" when X = 12 AND Y = 6 else
"100010011100" when X = 13 AND Y = 6 else
"100010001100" when X = 14 AND Y = 6 else
"101110101010" when X = 15 AND Y = 6 else
"111110010011" when X = 16 AND Y = 6 else
"111101000001" when X = 17 AND Y = 6 else
"101010001000" when X = 18 AND Y = 6 else
"000001001111" when X = 19 AND Y = 6 else
"001101001101" when X = 20 AND Y = 6 else
"111011100011" when X = 21 AND Y = 6 else
"111011110001" when X = 22 AND Y = 6 else
"110011010101" when X = 23 AND Y = 6 else
"000100101110" when X = 24 AND Y = 6 else
"000001101110" when X = 25 AND Y = 6 else
"110001110110" when X = 26 AND Y = 6 else
"111101000000" when X = 27 AND Y = 6 else
"111110010011" when X = 28 AND Y = 6 else
"101110101010" when X = 29 AND Y = 6 else
"100010001100" when X = 30 AND Y = 6 else
"100010011100" when X = 31 AND Y = 6 else
"111111110000" when X = 32 AND Y = 6 else
"100011001100" when X = 33 AND Y = 6 else
"001101000100" when X = 34 AND Y = 6 else
"000000000000" when X = 35 AND Y = 6 else
"001100110011" when X = 36 AND Y = 6 else
"010001010101" when X = 37 AND Y = 6 else
"011110101011" when X = 38 AND Y = 6 else
"111111110000" when X = 39 AND Y = 6 else
"111111110000" when X = 40 AND Y = 6 else
"111111110000" when X = 41 AND Y = 6 else
"111111110000" when X = 42 AND Y = 6 else
"111111110000" when X = 43 AND Y = 6 else
"111111110000" when X = 44 AND Y = 6 else
"111111110000" when X = 45 AND Y = 6 else
"111111110000" when X = 0 AND Y = 7 else
"111111110000" when X = 1 AND Y = 7 else
"111111110000" when X = 2 AND Y = 7 else
"111111110000" when X = 3 AND Y = 7 else
"111111110000" when X = 4 AND Y = 7 else
"111111110000" when X = 5 AND Y = 7 else
"001101010101" when X = 6 AND Y = 7 else
"001100110011" when X = 7 AND Y = 7 else
"001000100010" when X = 8 AND Y = 7 else
"000000000000" when X = 9 AND Y = 7 else
"000000000000" when X = 10 AND Y = 7 else
"010101000111" when X = 11 AND Y = 7 else
"100001011011" when X = 12 AND Y = 7 else
"100100111000" when X = 13 AND Y = 7 else
"110001010101" when X = 14 AND Y = 7 else
"111010000010" when X = 15 AND Y = 7 else
"111101110000" when X = 16 AND Y = 7 else
"110101000100" when X = 17 AND Y = 7 else
"010101111100" when X = 18 AND Y = 7 else
"000100111111" when X = 19 AND Y = 7 else
"100010011001" when X = 20 AND Y = 7 else
"111011100001" when X = 21 AND Y = 7 else
"111111110000" when X = 22 AND Y = 7 else
"111011100010" when X = 23 AND Y = 7 else
"011110001010" when X = 24 AND Y = 7 else
"000100111111" when X = 25 AND Y = 7 else
"011010001011" when X = 26 AND Y = 7 else
"110101010100" when X = 27 AND Y = 7 else
"111101110000" when X = 28 AND Y = 7 else
"111010000010" when X = 29 AND Y = 7 else
"110001010101" when X = 30 AND Y = 7 else
"100100111000" when X = 31 AND Y = 7 else
"100001011011" when X = 32 AND Y = 7 else
"011001000111" when X = 33 AND Y = 7 else
"000000000000" when X = 34 AND Y = 7 else
"000000000000" when X = 35 AND Y = 7 else
"001100110011" when X = 36 AND Y = 7 else
"001000100010" when X = 37 AND Y = 7 else
"010101110111" when X = 38 AND Y = 7 else
"111111110000" when X = 39 AND Y = 7 else
"111111110000" when X = 40 AND Y = 7 else
"111111110000" when X = 41 AND Y = 7 else
"111111110000" when X = 42 AND Y = 7 else
"111111110000" when X = 43 AND Y = 7 else
"111111110000" when X = 44 AND Y = 7 else
"111111110000" when X = 45 AND Y = 7 else
"111111110000" when X = 0 AND Y = 8 else
"111111110000" when X = 1 AND Y = 8 else
"111111110000" when X = 2 AND Y = 8 else
"111111110000" when X = 3 AND Y = 8 else
"111111110000" when X = 4 AND Y = 8 else
"111111110000" when X = 5 AND Y = 8 else
"001101010101" when X = 6 AND Y = 8 else
"000000000000" when X = 7 AND Y = 8 else
"000000000000" when X = 8 AND Y = 8 else
"000000000000" when X = 9 AND Y = 8 else
"011000110000" when X = 10 AND Y = 8 else
"110101110011" when X = 11 AND Y = 8 else
"110101100100" when X = 12 AND Y = 8 else
"111001110011" when X = 13 AND Y = 8 else
"111110010000" when X = 14 AND Y = 8 else
"111110010000" when X = 15 AND Y = 8 else
"111101110000" when X = 16 AND Y = 8 else
"101101110110" when X = 17 AND Y = 8 else
"000001101111" when X = 18 AND Y = 8 else
"001000111101" when X = 19 AND Y = 8 else
"110111010100" when X = 20 AND Y = 8 else
"111111100000" when X = 21 AND Y = 8 else
"111111100000" when X = 22 AND Y = 8 else
"111111100000" when X = 23 AND Y = 8 else
"101110110110" when X = 24 AND Y = 8 else
"000100011110" when X = 25 AND Y = 8 else
"000010001110" when X = 26 AND Y = 8 else
"101110000110" when X = 27 AND Y = 8 else
"111101110000" when X = 28 AND Y = 8 else
"111110010000" when X = 29 AND Y = 8 else
"111110010000" when X = 30 AND Y = 8 else
"111001110011" when X = 31 AND Y = 8 else
"110101100100" when X = 32 AND Y = 8 else
"110101110011" when X = 33 AND Y = 8 else
"011000110000" when X = 34 AND Y = 8 else
"000000000000" when X = 35 AND Y = 8 else
"000000000000" when X = 36 AND Y = 8 else
"000000000000" when X = 37 AND Y = 8 else
"010101110111" when X = 38 AND Y = 8 else
"111111110000" when X = 39 AND Y = 8 else
"111111110000" when X = 40 AND Y = 8 else
"111111110000" when X = 41 AND Y = 8 else
"111111110000" when X = 42 AND Y = 8 else
"111111110000" when X = 43 AND Y = 8 else
"111111110000" when X = 44 AND Y = 8 else
"111111110000" when X = 45 AND Y = 8 else
"111111110000" when X = 0 AND Y = 9 else
"111111110000" when X = 1 AND Y = 9 else
"111111110000" when X = 2 AND Y = 9 else
"111111110000" when X = 3 AND Y = 9 else
"111111110000" when X = 4 AND Y = 9 else
"111111110000" when X = 5 AND Y = 9 else
"001101010101" when X = 6 AND Y = 9 else
"000000000000" when X = 7 AND Y = 9 else
"000100000000" when X = 8 AND Y = 9 else
"011100110000" when X = 9 AND Y = 9 else
"111010000000" when X = 10 AND Y = 9 else
"111110000000" when X = 11 AND Y = 9 else
"111110000000" when X = 12 AND Y = 9 else
"111110010000" when X = 13 AND Y = 9 else
"111110010000" when X = 14 AND Y = 9 else
"111110010000" when X = 15 AND Y = 9 else
"110110010100" when X = 16 AND Y = 9 else
"010011001100" when X = 17 AND Y = 9 else
"001110001100" when X = 18 AND Y = 9 else
"101101110110" when X = 19 AND Y = 9 else
"111110010000" when X = 20 AND Y = 9 else
"111110010000" when X = 21 AND Y = 9 else
"111110010000" when X = 22 AND Y = 9 else
"111110010000" when X = 23 AND Y = 9 else
"111110010001" when X = 24 AND Y = 9 else
"100101101000" when X = 25 AND Y = 9 else
"001010011101" when X = 26 AND Y = 9 else
"010011001100" when X = 27 AND Y = 9 else
"110110010100" when X = 28 AND Y = 9 else
"111110010000" when X = 29 AND Y = 9 else
"111110010000" when X = 30 AND Y = 9 else
"111110010000" when X = 31 AND Y = 9 else
"111110000000" when X = 32 AND Y = 9 else
"111110000000" when X = 33 AND Y = 9 else
"111110000000" when X = 34 AND Y = 9 else
"011000110000" when X = 35 AND Y = 9 else
"000000000000" when X = 36 AND Y = 9 else
"000000000000" when X = 37 AND Y = 9 else
"010101110111" when X = 38 AND Y = 9 else
"111111110000" when X = 39 AND Y = 9 else
"111111110000" when X = 40 AND Y = 9 else
"111111110000" when X = 41 AND Y = 9 else
"111111110000" when X = 42 AND Y = 9 else
"111111110000" when X = 43 AND Y = 9 else
"111111110000" when X = 44 AND Y = 9 else
"111111110000" when X = 45 AND Y = 9 else
"111111110000" when X = 0 AND Y = 10 else
"111111110000" when X = 1 AND Y = 10 else
"111111110000" when X = 2 AND Y = 10 else
"111111110000" when X = 3 AND Y = 10 else
"111111110000" when X = 4 AND Y = 10 else
"111111110000" when X = 5 AND Y = 10 else
"001101000101" when X = 6 AND Y = 10 else
"000000000000" when X = 7 AND Y = 10 else
"100001000000" when X = 8 AND Y = 10 else
"111110000000" when X = 9 AND Y = 10 else
"111110000000" when X = 10 AND Y = 10 else
"111101000000" when X = 11 AND Y = 10 else
"111101010000" when X = 12 AND Y = 10 else
"111101100000" when X = 13 AND Y = 10 else
"111101100000" when X = 14 AND Y = 10 else
"111101100000" when X = 15 AND Y = 10 else
"111001100011" when X = 16 AND Y = 10 else
"100110001000" when X = 17 AND Y = 10 else
"110101110101" when X = 18 AND Y = 10 else
"111101100000" when X = 19 AND Y = 10 else
"111101100000" when X = 20 AND Y = 10 else
"111101100000" when X = 21 AND Y = 10 else
"111101100000" when X = 22 AND Y = 10 else
"111101100000" when X = 23 AND Y = 10 else
"111101100000" when X = 24 AND Y = 10 else
"111101100000" when X = 25 AND Y = 10 else
"101101110110" when X = 26 AND Y = 10 else
"100110001000" when X = 27 AND Y = 10 else
"111001100011" when X = 28 AND Y = 10 else
"111101100000" when X = 29 AND Y = 10 else
"111101100000" when X = 30 AND Y = 10 else
"111101100000" when X = 31 AND Y = 10 else
"111101010000" when X = 32 AND Y = 10 else
"111101000000" when X = 33 AND Y = 10 else
"111110000000" when X = 34 AND Y = 10 else
"111110000000" when X = 35 AND Y = 10 else
"011000110000" when X = 36 AND Y = 10 else
"000000000000" when X = 37 AND Y = 10 else
"010101110111" when X = 38 AND Y = 10 else
"111111110000" when X = 39 AND Y = 10 else
"111111110000" when X = 40 AND Y = 10 else
"111111110000" when X = 41 AND Y = 10 else
"111111110000" when X = 42 AND Y = 10 else
"111111110000" when X = 43 AND Y = 10 else
"111111110000" when X = 44 AND Y = 10 else
"111111110000" when X = 45 AND Y = 10 else
"111111110000" when X = 0 AND Y = 11 else
"111111110000" when X = 1 AND Y = 11 else
"111111110000" when X = 2 AND Y = 11 else
"111111110000" when X = 3 AND Y = 11 else
"111111110000" when X = 4 AND Y = 11 else
"101111001011" when X = 5 AND Y = 11 else
"101001100011" when X = 6 AND Y = 11 else
"100101010000" when X = 7 AND Y = 11 else
"111010000000" when X = 8 AND Y = 11 else
"111110000000" when X = 9 AND Y = 11 else
"111110000000" when X = 10 AND Y = 11 else
"111101000000" when X = 11 AND Y = 11 else
"110000000000" when X = 12 AND Y = 11 else
"101100000000" when X = 13 AND Y = 11 else
"101100000000" when X = 14 AND Y = 11 else
"101100000000" when X = 15 AND Y = 11 else
"101100000000" when X = 16 AND Y = 11 else
"101100000000" when X = 17 AND Y = 11 else
"101100000000" when X = 18 AND Y = 11 else
"101100000000" when X = 19 AND Y = 11 else
"101100000000" when X = 20 AND Y = 11 else
"101100000000" when X = 21 AND Y = 11 else
"101100000000" when X = 22 AND Y = 11 else
"101100000000" when X = 23 AND Y = 11 else
"101100000000" when X = 24 AND Y = 11 else
"101100000000" when X = 25 AND Y = 11 else
"101100000000" when X = 26 AND Y = 11 else
"101100000000" when X = 27 AND Y = 11 else
"101100000000" when X = 28 AND Y = 11 else
"101100000000" when X = 29 AND Y = 11 else
"101100000000" when X = 30 AND Y = 11 else
"101100000000" when X = 31 AND Y = 11 else
"110000000000" when X = 32 AND Y = 11 else
"111101000000" when X = 33 AND Y = 11 else
"111110000000" when X = 34 AND Y = 11 else
"111110000000" when X = 35 AND Y = 11 else
"111010000000" when X = 36 AND Y = 11 else
"100101010000" when X = 37 AND Y = 11 else
"101110000100" when X = 38 AND Y = 11 else
"101011001100" when X = 39 AND Y = 11 else
"111111110000" when X = 40 AND Y = 11 else
"111111110000" when X = 41 AND Y = 11 else
"111111110000" when X = 42 AND Y = 11 else
"111111110000" when X = 43 AND Y = 11 else
"111111110000" when X = 44 AND Y = 11 else
"111111110000" when X = 45 AND Y = 11 else
"111111110000" when X = 0 AND Y = 12 else
"111111110000" when X = 1 AND Y = 12 else
"010101110111" when X = 2 AND Y = 12 else
"001000110011" when X = 3 AND Y = 12 else
"001000110011" when X = 4 AND Y = 12 else
"001100100010" when X = 5 AND Y = 12 else
"010000100000" when X = 6 AND Y = 12 else
"010000100000" when X = 7 AND Y = 12 else
"001100100000" when X = 8 AND Y = 12 else
"011101000000" when X = 9 AND Y = 12 else
"111110000000" when X = 10 AND Y = 12 else
"111101000000" when X = 11 AND Y = 12 else
"101000000000" when X = 12 AND Y = 12 else
"100000000000" when X = 13 AND Y = 12 else
"100000000000" when X = 14 AND Y = 12 else
"100000000000" when X = 15 AND Y = 12 else
"100000000000" when X = 16 AND Y = 12 else
"100000000000" when X = 17 AND Y = 12 else
"100000000000" when X = 18 AND Y = 12 else
"100000000000" when X = 19 AND Y = 12 else
"100000000000" when X = 20 AND Y = 12 else
"100000000000" when X = 21 AND Y = 12 else
"100100000000" when X = 22 AND Y = 12 else
"100000000000" when X = 23 AND Y = 12 else
"100000000000" when X = 24 AND Y = 12 else
"100000000000" when X = 25 AND Y = 12 else
"100000000000" when X = 26 AND Y = 12 else
"100000000000" when X = 27 AND Y = 12 else
"100000000000" when X = 28 AND Y = 12 else
"100000000000" when X = 29 AND Y = 12 else
"100000000000" when X = 30 AND Y = 12 else
"100000000000" when X = 31 AND Y = 12 else
"101000000000" when X = 32 AND Y = 12 else
"111101000000" when X = 33 AND Y = 12 else
"111110000000" when X = 34 AND Y = 12 else
"011101000000" when X = 35 AND Y = 12 else
"001100100000" when X = 36 AND Y = 12 else
"010000100000" when X = 37 AND Y = 12 else
"010000100000" when X = 38 AND Y = 12 else
"001000110010" when X = 39 AND Y = 12 else
"001000110011" when X = 40 AND Y = 12 else
"001000110011" when X = 41 AND Y = 12 else
"011010001001" when X = 42 AND Y = 12 else
"111111110000" when X = 43 AND Y = 12 else
"111111110000" when X = 44 AND Y = 12 else
"111111110000" when X = 45 AND Y = 12 else
"111111110000" when X = 0 AND Y = 13 else
"011010011010" when X = 1 AND Y = 13 else
"000000010001" when X = 2 AND Y = 13 else
"000000000000" when X = 3 AND Y = 13 else
"000000000000" when X = 4 AND Y = 13 else
"000000000000" when X = 5 AND Y = 13 else
"000100010001" when X = 6 AND Y = 13 else
"000100010001" when X = 7 AND Y = 13 else
"000000000000" when X = 8 AND Y = 13 else
"000100000000" when X = 9 AND Y = 13 else
"100001010010" when X = 10 AND Y = 13 else
"111100110001" when X = 11 AND Y = 13 else
"101000000000" when X = 12 AND Y = 13 else
"100100000000" when X = 13 AND Y = 13 else
"100100000000" when X = 14 AND Y = 13 else
"100100000000" when X = 15 AND Y = 13 else
"100100000000" when X = 16 AND Y = 13 else
"100100000000" when X = 17 AND Y = 13 else
"100100000000" when X = 18 AND Y = 13 else
"100100000000" when X = 19 AND Y = 13 else
"100000000000" when X = 20 AND Y = 13 else
"101100000000" when X = 21 AND Y = 13 else
"111000000000" when X = 22 AND Y = 13 else
"101000000000" when X = 23 AND Y = 13 else
"100000000000" when X = 24 AND Y = 13 else
"100100000000" when X = 25 AND Y = 13 else
"100100000000" when X = 26 AND Y = 13 else
"100100000000" when X = 27 AND Y = 13 else
"100100000000" when X = 28 AND Y = 13 else
"100100000000" when X = 29 AND Y = 13 else
"100100000000" when X = 30 AND Y = 13 else
"100100000000" when X = 31 AND Y = 13 else
"101000000000" when X = 32 AND Y = 13 else
"111100110001" when X = 33 AND Y = 13 else
"100101010010" when X = 34 AND Y = 13 else
"000100000000" when X = 35 AND Y = 13 else
"000000000001" when X = 36 AND Y = 13 else
"000100010001" when X = 37 AND Y = 13 else
"000100010001" when X = 38 AND Y = 13 else
"000000000000" when X = 39 AND Y = 13 else
"000100000000" when X = 40 AND Y = 13 else
"000000000000" when X = 41 AND Y = 13 else
"000100100010" when X = 42 AND Y = 13 else
"011110101011" when X = 43 AND Y = 13 else
"111111110000" when X = 44 AND Y = 13 else
"111111110000" when X = 45 AND Y = 13 else
"111111110000" when X = 0 AND Y = 14 else
"010101111000" when X = 1 AND Y = 14 else
"000000000000" when X = 2 AND Y = 14 else
"010001000100" when X = 3 AND Y = 14 else
"010001000100" when X = 4 AND Y = 14 else
"001000100010" when X = 5 AND Y = 14 else
"011001100110" when X = 6 AND Y = 14 else
"011001100110" when X = 7 AND Y = 14 else
"010001000100" when X = 8 AND Y = 14 else
"000000000000" when X = 9 AND Y = 14 else
"000100010111" when X = 10 AND Y = 14 else
"101000100110" when X = 11 AND Y = 14 else
"100000010011" when X = 12 AND Y = 14 else
"011000000100" when X = 13 AND Y = 14 else
"011000000100" when X = 14 AND Y = 14 else
"011000000100" when X = 15 AND Y = 14 else
"011000000100" when X = 16 AND Y = 14 else
"011000000100" when X = 17 AND Y = 14 else
"011000000100" when X = 18 AND Y = 14 else
"011000000100" when X = 19 AND Y = 14 else
"011100000011" when X = 20 AND Y = 14 else
"110000000000" when X = 21 AND Y = 14 else
"111100000000" when X = 22 AND Y = 14 else
"101100000001" when X = 23 AND Y = 14 else
"011000000100" when X = 24 AND Y = 14 else
"011000000100" when X = 25 AND Y = 14 else
"011000000100" when X = 26 AND Y = 14 else
"011000000100" when X = 27 AND Y = 14 else
"011000000100" when X = 28 AND Y = 14 else
"011000000100" when X = 29 AND Y = 14 else
"011000000100" when X = 30 AND Y = 14 else
"011000000100" when X = 31 AND Y = 14 else
"100000010011" when X = 32 AND Y = 14 else
"101000100110" when X = 33 AND Y = 14 else
"000100010111" when X = 34 AND Y = 14 else
"000000000000" when X = 35 AND Y = 14 else
"010101010101" when X = 36 AND Y = 14 else
"011001100110" when X = 37 AND Y = 14 else
"011001100110" when X = 38 AND Y = 14 else
"001000100010" when X = 39 AND Y = 14 else
"010101010101" when X = 40 AND Y = 14 else
"001100110011" when X = 41 AND Y = 14 else
"000000000000" when X = 42 AND Y = 14 else
"011110101010" when X = 43 AND Y = 14 else
"111111110000" when X = 44 AND Y = 14 else
"111111110000" when X = 45 AND Y = 14 else
"111111110000" when X = 0 AND Y = 15 else
"010101111000" when X = 1 AND Y = 15 else
"000000000000" when X = 2 AND Y = 15 else
"000000000000" when X = 3 AND Y = 15 else
"000000000000" when X = 4 AND Y = 15 else
"000000000000" when X = 5 AND Y = 15 else
"000000000000" when X = 6 AND Y = 15 else
"000000000000" when X = 7 AND Y = 15 else
"000000000000" when X = 8 AND Y = 15 else
"000000000000" when X = 9 AND Y = 15 else
"000000000111" when X = 10 AND Y = 15 else
"100100010111" when X = 11 AND Y = 15 else
"001100011100" when X = 12 AND Y = 15 else
"000100101110" when X = 13 AND Y = 15 else
"000001001100" when X = 14 AND Y = 15 else
"000001001100" when X = 15 AND Y = 15 else
"000101001100" when X = 16 AND Y = 15 else
"001100011100" when X = 17 AND Y = 15 else
"001000111100" when X = 18 AND Y = 15 else
"001000101101" when X = 19 AND Y = 15 else
"011000011010" when X = 20 AND Y = 15 else
"111100000001" when X = 21 AND Y = 15 else
"111100000000" when X = 22 AND Y = 15 else
"111000000010" when X = 23 AND Y = 15 else
"010000011011" when X = 24 AND Y = 15 else
"001000101100" when X = 25 AND Y = 15 else
"001000101100" when X = 26 AND Y = 15 else
"001100011100" when X = 27 AND Y = 15 else
"000101001100" when X = 28 AND Y = 15 else
"000001001100" when X = 29 AND Y = 15 else
"000101001100" when X = 30 AND Y = 15 else
"000100101110" when X = 31 AND Y = 15 else
"001100011101" when X = 32 AND Y = 15 else
"100100010111" when X = 33 AND Y = 15 else
"000000000111" when X = 34 AND Y = 15 else
"000000000000" when X = 35 AND Y = 15 else
"000000000000" when X = 36 AND Y = 15 else
"000000000000" when X = 37 AND Y = 15 else
"000000000000" when X = 38 AND Y = 15 else
"000000000000" when X = 39 AND Y = 15 else
"000000000000" when X = 40 AND Y = 15 else
"000000000000" when X = 41 AND Y = 15 else
"000000000000" when X = 42 AND Y = 15 else
"011110101010" when X = 43 AND Y = 15 else
"111111110000" when X = 44 AND Y = 15 else
"111111110000" when X = 45 AND Y = 15 else
"111111110000" when X = 0 AND Y = 16 else
"010101111000" when X = 1 AND Y = 16 else
"000000000000" when X = 2 AND Y = 16 else
"000000000000" when X = 3 AND Y = 16 else
"000000000000" when X = 4 AND Y = 16 else
"000000000000" when X = 5 AND Y = 16 else
"000000000000" when X = 6 AND Y = 16 else
"000000000000" when X = 7 AND Y = 16 else
"000000000000" when X = 8 AND Y = 16 else
"000000000000" when X = 9 AND Y = 16 else
"001000000110" when X = 10 AND Y = 16 else
"010100011011" when X = 11 AND Y = 16 else
"000100001111" when X = 12 AND Y = 16 else
"000001001101" when X = 13 AND Y = 16 else
"000010011000" when X = 14 AND Y = 16 else
"000110001000" when X = 15 AND Y = 16 else
"010101001001" when X = 16 AND Y = 16 else
"011100011001" when X = 17 AND Y = 16 else
"010101011001" when X = 18 AND Y = 16 else
"010100111001" when X = 19 AND Y = 16 else
"100100001000" when X = 20 AND Y = 16 else
"111100000000" when X = 21 AND Y = 16 else
"111100000000" when X = 22 AND Y = 16 else
"111000000010" when X = 23 AND Y = 16 else
"100000001000" when X = 24 AND Y = 16 else
"010101001001" when X = 25 AND Y = 16 else
"010101001001" when X = 26 AND Y = 16 else
"011100001001" when X = 27 AND Y = 16 else
"010101001001" when X = 28 AND Y = 16 else
"000110001000" when X = 29 AND Y = 16 else
"000010011000" when X = 30 AND Y = 16 else
"000001001101" when X = 31 AND Y = 16 else
"000100001111" when X = 32 AND Y = 16 else
"010100011011" when X = 33 AND Y = 16 else
"001000000110" when X = 34 AND Y = 16 else
"000000000000" when X = 35 AND Y = 16 else
"000000000000" when X = 36 AND Y = 16 else
"000000000000" when X = 37 AND Y = 16 else
"000000000000" when X = 38 AND Y = 16 else
"000000000000" when X = 39 AND Y = 16 else
"000000000000" when X = 40 AND Y = 16 else
"000000000000" when X = 41 AND Y = 16 else
"000000000000" when X = 42 AND Y = 16 else
"011110101010" when X = 43 AND Y = 16 else
"111111110000" when X = 44 AND Y = 16 else
"111111110000" when X = 45 AND Y = 16 else
"111111110000" when X = 0 AND Y = 17 else
"010101111000" when X = 1 AND Y = 17 else
"000000000000" when X = 2 AND Y = 17 else
"000000000000" when X = 3 AND Y = 17 else
"000000000000" when X = 4 AND Y = 17 else
"000000000000" when X = 5 AND Y = 17 else
"000000000000" when X = 6 AND Y = 17 else
"000000000000" when X = 7 AND Y = 17 else
"000000000000" when X = 8 AND Y = 17 else
"000000000000" when X = 9 AND Y = 17 else
"001100000100" when X = 10 AND Y = 17 else
"010100001011" when X = 11 AND Y = 17 else
"001000101101" when X = 12 AND Y = 17 else
"001001101010" when X = 13 AND Y = 17 else
"001010001001" when X = 14 AND Y = 17 else
"001101111001" when X = 15 AND Y = 17 else
"011000101001" when X = 16 AND Y = 17 else
"011100001001" when X = 17 AND Y = 17 else
"010001011001" when X = 18 AND Y = 17 else
"011001001001" when X = 19 AND Y = 17 else
"100100101000" when X = 20 AND Y = 17 else
"111100100010" when X = 21 AND Y = 17 else
"111100100001" when X = 22 AND Y = 17 else
"111000100011" when X = 23 AND Y = 17 else
"100000101001" when X = 24 AND Y = 17 else
"010101011001" when X = 25 AND Y = 17 else
"010101001001" when X = 26 AND Y = 17 else
"011100001001" when X = 27 AND Y = 17 else
"011000101001" when X = 28 AND Y = 17 else
"001101111001" when X = 29 AND Y = 17 else
"001010001001" when X = 30 AND Y = 17 else
"001001101010" when X = 31 AND Y = 17 else
"001000101101" when X = 32 AND Y = 17 else
"010100001011" when X = 33 AND Y = 17 else
"001100000100" when X = 34 AND Y = 17 else
"000000000000" when X = 35 AND Y = 17 else
"000000000000" when X = 36 AND Y = 17 else
"000000000000" when X = 37 AND Y = 17 else
"000000000000" when X = 38 AND Y = 17 else
"000000000000" when X = 39 AND Y = 17 else
"000000000000" when X = 40 AND Y = 17 else
"000000000000" when X = 41 AND Y = 17 else
"000000000000" when X = 42 AND Y = 17 else
"011110101010" when X = 43 AND Y = 17 else
"111111110000" when X = 44 AND Y = 17 else
"111111110000" when X = 45 AND Y = 17 else
"111111110000" when X = 0 AND Y = 18 else
"011010001001" when X = 1 AND Y = 18 else
"000000000000" when X = 2 AND Y = 18 else
"000000000000" when X = 3 AND Y = 18 else
"000000000000" when X = 4 AND Y = 18 else
"000000000000" when X = 5 AND Y = 18 else
"000000000000" when X = 6 AND Y = 18 else
"000000000000" when X = 7 AND Y = 18 else
"000000000000" when X = 8 AND Y = 18 else
"000000000000" when X = 9 AND Y = 18 else
"001100000100" when X = 10 AND Y = 18 else
"011100001001" when X = 11 AND Y = 18 else
"011000011010" when X = 12 AND Y = 18 else
"011000101001" when X = 13 AND Y = 18 else
"011000101001" when X = 14 AND Y = 18 else
"011000011001" when X = 15 AND Y = 18 else
"011000011001" when X = 16 AND Y = 18 else
"011100001001" when X = 17 AND Y = 18 else
"010101011001" when X = 18 AND Y = 18 else
"011110011001" when X = 19 AND Y = 18 else
"101010001001" when X = 20 AND Y = 18 else
"101010011000" when X = 21 AND Y = 18 else
"101010011000" when X = 22 AND Y = 18 else
"101010001001" when X = 23 AND Y = 18 else
"100110001001" when X = 24 AND Y = 18 else
"011010001001" when X = 25 AND Y = 18 else
"010101001001" when X = 26 AND Y = 18 else
"011100001001" when X = 27 AND Y = 18 else
"011000011001" when X = 28 AND Y = 18 else
"011000011001" when X = 29 AND Y = 18 else
"011000101001" when X = 30 AND Y = 18 else
"011000101001" when X = 31 AND Y = 18 else
"011000011010" when X = 32 AND Y = 18 else
"011100001001" when X = 33 AND Y = 18 else
"001100000100" when X = 34 AND Y = 18 else
"000000000000" when X = 35 AND Y = 18 else
"000000000000" when X = 36 AND Y = 18 else
"000000000000" when X = 37 AND Y = 18 else
"000000000000" when X = 38 AND Y = 18 else
"000000000000" when X = 39 AND Y = 18 else
"000000000000" when X = 40 AND Y = 18 else
"000000000000" when X = 41 AND Y = 18 else
"000100010001" when X = 42 AND Y = 18 else
"011110101011" when X = 43 AND Y = 18 else
"111111110000" when X = 44 AND Y = 18 else
"111111110000" when X = 45 AND Y = 18 else
"111111110000" when X = 0 AND Y = 19 else
"100110111100" when X = 1 AND Y = 19 else
"001100110011" when X = 2 AND Y = 19 else
"000000000000" when X = 3 AND Y = 19 else
"000000000000" when X = 4 AND Y = 19 else
"000000000000" when X = 5 AND Y = 19 else
"000000000000" when X = 6 AND Y = 19 else
"000000000000" when X = 7 AND Y = 19 else
"000000000000" when X = 8 AND Y = 19 else
"000000000000" when X = 9 AND Y = 19 else
"001100000100" when X = 10 AND Y = 19 else
"011000001010" when X = 11 AND Y = 19 else
"010000011011" when X = 12 AND Y = 19 else
"010101001001" when X = 13 AND Y = 19 else
"010101001001" when X = 14 AND Y = 19 else
"010101001001" when X = 15 AND Y = 19 else
"011000011001" when X = 16 AND Y = 19 else
"011100001001" when X = 17 AND Y = 19 else
"010101011001" when X = 18 AND Y = 19 else
"011110011001" when X = 19 AND Y = 19 else
"011110011001" when X = 20 AND Y = 19 else
"011010011001" when X = 21 AND Y = 19 else
"011010011001" when X = 22 AND Y = 19 else
"011010011001" when X = 23 AND Y = 19 else
"011110011001" when X = 24 AND Y = 19 else
"011010011001" when X = 25 AND Y = 19 else
"010101001001" when X = 26 AND Y = 19 else
"011100001001" when X = 27 AND Y = 19 else
"011000011001" when X = 28 AND Y = 19 else
"010101001001" when X = 29 AND Y = 19 else
"010101001001" when X = 30 AND Y = 19 else
"010101001001" when X = 31 AND Y = 19 else
"010000011011" when X = 32 AND Y = 19 else
"011000001010" when X = 33 AND Y = 19 else
"001100000100" when X = 34 AND Y = 19 else
"000000000000" when X = 35 AND Y = 19 else
"000000000000" when X = 36 AND Y = 19 else
"000000000000" when X = 37 AND Y = 19 else
"000000000000" when X = 38 AND Y = 19 else
"000000000000" when X = 39 AND Y = 19 else
"000000000000" when X = 40 AND Y = 19 else
"000000000000" when X = 41 AND Y = 19 else
"010101010101" when X = 42 AND Y = 19 else
"111011010101" when X = 43 AND Y = 19 else
"111111110000" when X = 44 AND Y = 19 else
"111111110000" when X = 45 AND Y = 19 else
"111111110000" when X = 0 AND Y = 20 else
"100110111100" when X = 1 AND Y = 20 else
"001100110011" when X = 2 AND Y = 20 else
"000000000000" when X = 3 AND Y = 20 else
"000000000000" when X = 4 AND Y = 20 else
"000000000000" when X = 5 AND Y = 20 else
"000000000000" when X = 6 AND Y = 20 else
"000000000000" when X = 7 AND Y = 20 else
"000000000000" when X = 8 AND Y = 20 else
"000000000000" when X = 9 AND Y = 20 else
"001100000101" when X = 10 AND Y = 20 else
"010000011100" when X = 11 AND Y = 20 else
"000101011011" when X = 12 AND Y = 20 else
"000010001001" when X = 13 AND Y = 20 else
"000010011000" when X = 14 AND Y = 20 else
"000110001001" when X = 15 AND Y = 20 else
"011000101001" when X = 16 AND Y = 20 else
"011000001001" when X = 17 AND Y = 20 else
"010101011001" when X = 18 AND Y = 20 else
"011010011001" when X = 19 AND Y = 20 else
"001010011001" when X = 20 AND Y = 20 else
"000001111010" when X = 21 AND Y = 20 else
"000001001101" when X = 22 AND Y = 20 else
"000001111010" when X = 23 AND Y = 20 else
"010010011001" when X = 24 AND Y = 20 else
"011010011001" when X = 25 AND Y = 20 else
"010101001001" when X = 26 AND Y = 20 else
"011000001001" when X = 27 AND Y = 20 else
"011000101001" when X = 28 AND Y = 20 else
"000110001001" when X = 29 AND Y = 20 else
"000010011000" when X = 30 AND Y = 20 else
"000010001001" when X = 31 AND Y = 20 else
"000101011011" when X = 32 AND Y = 20 else
"010000011100" when X = 33 AND Y = 20 else
"001100000101" when X = 34 AND Y = 20 else
"000000000000" when X = 35 AND Y = 20 else
"000000000000" when X = 36 AND Y = 20 else
"000000000000" when X = 37 AND Y = 20 else
"000000000000" when X = 38 AND Y = 20 else
"000000000000" when X = 39 AND Y = 20 else
"000000000000" when X = 40 AND Y = 20 else
"000000000000" when X = 41 AND Y = 20 else
"010101010101" when X = 42 AND Y = 20 else
"111011010101" when X = 43 AND Y = 20 else
"111111110000" when X = 44 AND Y = 20 else
"111111110000" when X = 45 AND Y = 20 else
"111111110000" when X = 0 AND Y = 21 else
"011010001001" when X = 1 AND Y = 21 else
"000000000000" when X = 2 AND Y = 21 else
"000000000000" when X = 3 AND Y = 21 else
"000000000000" when X = 4 AND Y = 21 else
"000000000000" when X = 5 AND Y = 21 else
"000000000000" when X = 6 AND Y = 21 else
"000000000000" when X = 7 AND Y = 21 else
"000000000000" when X = 8 AND Y = 21 else
"000000000000" when X = 9 AND Y = 21 else
"000100010111" when X = 10 AND Y = 21 else
"000100011111" when X = 11 AND Y = 21 else
"000001111010" when X = 12 AND Y = 21 else
"000010011000" when X = 13 AND Y = 21 else
"000010001001" when X = 14 AND Y = 21 else
"000001001101" when X = 15 AND Y = 21 else
"001000001110" when X = 16 AND Y = 21 else
"001100001101" when X = 17 AND Y = 21 else
"010001011001" when X = 18 AND Y = 21 else
"011010011001" when X = 19 AND Y = 21 else
"001010011001" when X = 20 AND Y = 21 else
"000001101011" when X = 21 AND Y = 21 else
"000100101111" when X = 22 AND Y = 21 else
"000001111010" when X = 23 AND Y = 21 else
"010010011001" when X = 24 AND Y = 21 else
"011010011001" when X = 25 AND Y = 21 else
"010101001001" when X = 26 AND Y = 21 else
"001100001101" when X = 27 AND Y = 21 else
"001000001110" when X = 28 AND Y = 21 else
"000001001101" when X = 29 AND Y = 21 else
"000010001001" when X = 30 AND Y = 21 else
"000010011000" when X = 31 AND Y = 21 else
"000001111010" when X = 32 AND Y = 21 else
"000100011111" when X = 33 AND Y = 21 else
"000100010111" when X = 34 AND Y = 21 else
"000000000000" when X = 35 AND Y = 21 else
"000000000000" when X = 36 AND Y = 21 else
"000000000000" when X = 37 AND Y = 21 else
"000000000000" when X = 38 AND Y = 21 else
"000000000000" when X = 39 AND Y = 21 else
"000000000000" when X = 40 AND Y = 21 else
"000000000000" when X = 41 AND Y = 21 else
"000100010001" when X = 42 AND Y = 21 else
"011110101011" when X = 43 AND Y = 21 else
"111111110000" when X = 44 AND Y = 21 else
"111111110000" when X = 45 AND Y = 21 else
"111111110000" when X = 0 AND Y = 22 else
"010101111000" when X = 1 AND Y = 22 else
"000000000000" when X = 2 AND Y = 22 else
"000000000000" when X = 3 AND Y = 22 else
"000000000000" when X = 4 AND Y = 22 else
"000000000000" when X = 5 AND Y = 22 else
"000000000000" when X = 6 AND Y = 22 else
"000000000000" when X = 7 AND Y = 22 else
"000000000000" when X = 8 AND Y = 22 else
"000000000000" when X = 9 AND Y = 22 else
"010001010111" when X = 10 AND Y = 22 else
"010001111111" when X = 11 AND Y = 22 else
"000000111110" when X = 12 AND Y = 22 else
"000001111010" when X = 13 AND Y = 22 else
"000001011100" when X = 14 AND Y = 22 else
"000100001111" when X = 15 AND Y = 22 else
"000100001111" when X = 16 AND Y = 22 else
"000100001111" when X = 17 AND Y = 22 else
"000101011011" when X = 18 AND Y = 22 else
"011110011001" when X = 19 AND Y = 22 else
"001010011001" when X = 20 AND Y = 22 else
"000010001001" when X = 21 AND Y = 22 else
"000010001001" when X = 22 AND Y = 22 else
"000010001001" when X = 23 AND Y = 22 else
"010010011001" when X = 24 AND Y = 22 else
"011010011001" when X = 25 AND Y = 22 else
"000101001100" when X = 26 AND Y = 22 else
"000100001111" when X = 27 AND Y = 22 else
"000100001111" when X = 28 AND Y = 22 else
"000100001111" when X = 29 AND Y = 22 else
"000001011100" when X = 30 AND Y = 22 else
"000001111010" when X = 31 AND Y = 22 else
"000000111110" when X = 32 AND Y = 22 else
"010001111111" when X = 33 AND Y = 22 else
"010001100111" when X = 34 AND Y = 22 else
"000000000000" when X = 35 AND Y = 22 else
"000000000000" when X = 36 AND Y = 22 else
"000000000000" when X = 37 AND Y = 22 else
"000000000000" when X = 38 AND Y = 22 else
"000000000000" when X = 39 AND Y = 22 else
"000000000000" when X = 40 AND Y = 22 else
"000000000000" when X = 41 AND Y = 22 else
"000000000000" when X = 42 AND Y = 22 else
"011110101010" when X = 43 AND Y = 22 else
"111111110000" when X = 44 AND Y = 22 else
"111111110000" when X = 45 AND Y = 22 else
"111111110000" when X = 0 AND Y = 23 else
"010101111000" when X = 1 AND Y = 23 else
"000000000000" when X = 2 AND Y = 23 else
"000000000000" when X = 3 AND Y = 23 else
"000000000000" when X = 4 AND Y = 23 else
"000000000000" when X = 5 AND Y = 23 else
"000000000000" when X = 6 AND Y = 23 else
"000000000000" when X = 7 AND Y = 23 else
"000000000000" when X = 8 AND Y = 23 else
"000000000000" when X = 9 AND Y = 23 else
"010001100111" when X = 10 AND Y = 23 else
"111111110000" when X = 11 AND Y = 23 else
"010001101111" when X = 12 AND Y = 23 else
"000000111110" when X = 13 AND Y = 23 else
"000000111110" when X = 14 AND Y = 23 else
"000100001111" when X = 15 AND Y = 23 else
"000100001111" when X = 16 AND Y = 23 else
"000100001111" when X = 17 AND Y = 23 else
"000001011100" when X = 18 AND Y = 23 else
"011110011001" when X = 19 AND Y = 23 else
"011010011001" when X = 20 AND Y = 23 else
"010110011001" when X = 21 AND Y = 23 else
"010110011001" when X = 22 AND Y = 23 else
"010110011001" when X = 23 AND Y = 23 else
"011010011001" when X = 24 AND Y = 23 else
"011010011001" when X = 25 AND Y = 23 else
"000001001101" when X = 26 AND Y = 23 else
"000100001111" when X = 27 AND Y = 23 else
"000100001111" when X = 28 AND Y = 23 else
"000100001111" when X = 29 AND Y = 23 else
"000000111110" when X = 30 AND Y = 23 else
"000000111110" when X = 31 AND Y = 23 else
"001101101111" when X = 32 AND Y = 23 else
"111111110000" when X = 33 AND Y = 23 else
"010001100111" when X = 34 AND Y = 23 else
"000000000000" when X = 35 AND Y = 23 else
"000000000000" when X = 36 AND Y = 23 else
"000000000000" when X = 37 AND Y = 23 else
"000000000000" when X = 38 AND Y = 23 else
"000000000000" when X = 39 AND Y = 23 else
"000000000000" when X = 40 AND Y = 23 else
"000000000000" when X = 41 AND Y = 23 else
"000000000000" when X = 42 AND Y = 23 else
"011110101010" when X = 43 AND Y = 23 else
"111111110000" when X = 44 AND Y = 23 else
"111111110000" when X = 45 AND Y = 23 else
"111111110000" when X = 0 AND Y = 24 else
"010110001000" when X = 1 AND Y = 24 else
"000000000000" when X = 2 AND Y = 24 else
"000000000000" when X = 3 AND Y = 24 else
"000000000000" when X = 4 AND Y = 24 else
"000000000000" when X = 5 AND Y = 24 else
"000000000000" when X = 6 AND Y = 24 else
"000000000000" when X = 7 AND Y = 24 else
"000000000000" when X = 8 AND Y = 24 else
"000000000000" when X = 9 AND Y = 24 else
"010001100111" when X = 10 AND Y = 24 else
"111111110000" when X = 11 AND Y = 24 else
"111111110000" when X = 12 AND Y = 24 else
"010110011111" when X = 13 AND Y = 24 else
"010110001111" when X = 14 AND Y = 24 else
"001000111111" when X = 15 AND Y = 24 else
"000100001111" when X = 16 AND Y = 24 else
"001001001111" when X = 17 AND Y = 24 else
"011010101101" when X = 18 AND Y = 24 else
"100011001100" when X = 19 AND Y = 24 else
"100111001100" when X = 20 AND Y = 24 else
"100111001100" when X = 21 AND Y = 24 else
"100111001100" when X = 22 AND Y = 24 else
"100111001100" when X = 23 AND Y = 24 else
"100111001100" when X = 24 AND Y = 24 else
"100010111100" when X = 25 AND Y = 24 else
"010110011110" when X = 26 AND Y = 24 else
"001001001111" when X = 27 AND Y = 24 else
"000100001111" when X = 28 AND Y = 24 else
"001000111111" when X = 29 AND Y = 24 else
"010110001111" when X = 30 AND Y = 24 else
"010110011111" when X = 31 AND Y = 24 else
"111111110000" when X = 32 AND Y = 24 else
"111111110000" when X = 33 AND Y = 24 else
"010001110111" when X = 34 AND Y = 24 else
"000000000000" when X = 35 AND Y = 24 else
"000000000000" when X = 36 AND Y = 24 else
"000000000000" when X = 37 AND Y = 24 else
"000000000000" when X = 38 AND Y = 24 else
"000000000000" when X = 39 AND Y = 24 else
"000000000000" when X = 40 AND Y = 24 else
"000000000000" when X = 41 AND Y = 24 else
"000000000000" when X = 42 AND Y = 24 else
"011110101010" when X = 43 AND Y = 24 else
"111111110000" when X = 44 AND Y = 24 else
"111111110000" when X = 45 AND Y = 24 else
"111111110000" when X = 0 AND Y = 25 else
"100011001101" when X = 1 AND Y = 25 else
"001101010101" when X = 2 AND Y = 25 else
"000100010001" when X = 3 AND Y = 25 else
"000100010001" when X = 4 AND Y = 25 else
"000100010001" when X = 5 AND Y = 25 else
"000100010001" when X = 6 AND Y = 25 else
"000100010001" when X = 7 AND Y = 25 else
"000100010001" when X = 8 AND Y = 25 else
"001101000100" when X = 9 AND Y = 25 else
"100010111100" when X = 10 AND Y = 25 else
"111111110000" when X = 11 AND Y = 25 else
"111111110000" when X = 12 AND Y = 25 else
"111111110000" when X = 13 AND Y = 25 else
"111111110000" when X = 14 AND Y = 25 else
"011110111110" when X = 15 AND Y = 25 else
"011010101111" when X = 16 AND Y = 25 else
"100010111110" when X = 17 AND Y = 25 else
"111111110000" when X = 18 AND Y = 25 else
"111111110000" when X = 19 AND Y = 25 else
"111111110000" when X = 20 AND Y = 25 else
"111111110000" when X = 21 AND Y = 25 else
"111111110000" when X = 22 AND Y = 25 else
"111111110000" when X = 23 AND Y = 25 else
"111111110000" when X = 24 AND Y = 25 else
"111111110000" when X = 25 AND Y = 25 else
"111111110000" when X = 26 AND Y = 25 else
"100010111110" when X = 27 AND Y = 25 else
"011010101111" when X = 28 AND Y = 25 else
"011110111110" when X = 29 AND Y = 25 else
"111111110000" when X = 30 AND Y = 25 else
"111111110000" when X = 31 AND Y = 25 else
"111111110000" when X = 32 AND Y = 25 else
"111111110000" when X = 33 AND Y = 25 else
"100010111100" when X = 34 AND Y = 25 else
"001101000100" when X = 35 AND Y = 25 else
"000100010001" when X = 36 AND Y = 25 else
"000100010001" when X = 37 AND Y = 25 else
"000100010001" when X = 38 AND Y = 25 else
"000100010001" when X = 39 AND Y = 25 else
"000100010001" when X = 40 AND Y = 25 else
"000100010001" when X = 41 AND Y = 25 else
"010001100111" when X = 42 AND Y = 25 else
"111111110000" when X = 43 AND Y = 25 else
"111111110000" when X = 44 AND Y = 25 else
"111111110000" when X = 45 AND Y = 25 else
"111111110000" when X = 0 AND Y = 26 else
"111111110000" when X = 1 AND Y = 26 else
"111111110000" when X = 2 AND Y = 26 else
"100010111100" when X = 3 AND Y = 26 else
"100010111100" when X = 4 AND Y = 26 else
"100010111100" when X = 5 AND Y = 26 else
"100010111100" when X = 6 AND Y = 26 else
"100010111100" when X = 7 AND Y = 26 else
"100010111100" when X = 8 AND Y = 26 else
"111011010100" when X = 9 AND Y = 26 else
"111111110000" when X = 10 AND Y = 26 else
"111111110000" when X = 11 AND Y = 26 else
"111111110000" when X = 12 AND Y = 26 else
"111111110000" when X = 13 AND Y = 26 else
"111111110000" when X = 14 AND Y = 26 else
"111111110000" when X = 15 AND Y = 26 else
"111111110000" when X = 16 AND Y = 26 else
"111111110000" when X = 17 AND Y = 26 else
"111111110000" when X = 18 AND Y = 26 else
"111111110000" when X = 19 AND Y = 26 else
"111111110000" when X = 20 AND Y = 26 else
"111111110000" when X = 21 AND Y = 26 else
"111111110000" when X = 22 AND Y = 26 else
"111111110000" when X = 23 AND Y = 26 else
"111111110000" when X = 24 AND Y = 26 else
"111111110000" when X = 25 AND Y = 26 else
"111111110000" when X = 26 AND Y = 26 else
"111111110000" when X = 27 AND Y = 26 else
"111111110000" when X = 28 AND Y = 26 else
"111111110000" when X = 29 AND Y = 26 else
"111111110000" when X = 30 AND Y = 26 else
"111111110000" when X = 31 AND Y = 26 else
"111111110000" when X = 32 AND Y = 26 else
"111111110000" when X = 33 AND Y = 26 else
"111111110000" when X = 34 AND Y = 26 else
"111011010100" when X = 35 AND Y = 26 else
"100010111100" when X = 36 AND Y = 26 else
"100010111100" when X = 37 AND Y = 26 else
"100010111100" when X = 38 AND Y = 26 else
"100010111100" when X = 39 AND Y = 26 else
"100010111100" when X = 40 AND Y = 26 else
"100010111100" when X = 41 AND Y = 26 else
"111111110000" when X = 42 AND Y = 26 else
"111111110000" when X = 43 AND Y = 26 else
"111111110000" when X = 44 AND Y = 26 else
"111111110000" when X = 45 AND Y = 26 else
"111111110000" when X = 0 AND Y = 27 else
"111111110000" when X = 1 AND Y = 27 else
"111111110000" when X = 2 AND Y = 27 else
"111111110000" when X = 3 AND Y = 27 else
"111111110000" when X = 4 AND Y = 27 else
"111111110000" when X = 5 AND Y = 27 else
"111111110000" when X = 6 AND Y = 27 else
"111111110000" when X = 7 AND Y = 27 else
"111111110000" when X = 8 AND Y = 27 else
"111111110000" when X = 9 AND Y = 27 else
"111111110000" when X = 10 AND Y = 27 else
"111111110000" when X = 11 AND Y = 27 else
"111111110000" when X = 12 AND Y = 27 else
"111111110000" when X = 13 AND Y = 27 else
"111111110000" when X = 14 AND Y = 27 else
"111111110000" when X = 15 AND Y = 27 else
"111111110000" when X = 16 AND Y = 27 else
"111111110000" when X = 17 AND Y = 27 else
"111111110000" when X = 18 AND Y = 27 else
"111111110000" when X = 19 AND Y = 27 else
"111111110000" when X = 20 AND Y = 27 else
"111111110000" when X = 21 AND Y = 27 else
"111111110000" when X = 22 AND Y = 27 else
"111111110000" when X = 23 AND Y = 27 else
"111111110000" when X = 24 AND Y = 27 else
"111111110000" when X = 25 AND Y = 27 else
"111111110000" when X = 26 AND Y = 27 else
"111111110000" when X = 27 AND Y = 27 else
"111111110000" when X = 28 AND Y = 27 else
"111111110000" when X = 29 AND Y = 27 else
"111111110000" when X = 30 AND Y = 27 else
"111111110000" when X = 31 AND Y = 27 else
"111111110000" when X = 32 AND Y = 27 else
"111111110000" when X = 33 AND Y = 27 else
"111111110000" when X = 34 AND Y = 27 else
"111111110000" when X = 35 AND Y = 27 else
"111111110000" when X = 36 AND Y = 27 else
"111111110000" when X = 37 AND Y = 27 else
"111111110000" when X = 38 AND Y = 27 else
"111111110000" when X = 39 AND Y = 27 else
"111111110000" when X = 40 AND Y = 27 else
"111111110000" when X = 41 AND Y = 27 else
"111111110000" when X = 42 AND Y = 27 else
"111111110000" when X = 43 AND Y = 27 else
"111111110000" when X = 44 AND Y = 27 else
"111111110000" when X = 45 AND Y = 27 else
"111111110000" when X = 0 AND Y = 28 else
"111111110000" when X = 1 AND Y = 28 else
"111111110000" when X = 2 AND Y = 28 else
"111111110000" when X = 3 AND Y = 28 else
"111111110000" when X = 4 AND Y = 28 else
"111111110000" when X = 5 AND Y = 28 else
"111111110000" when X = 6 AND Y = 28 else
"111111110000" when X = 7 AND Y = 28 else
"111111110000" when X = 8 AND Y = 28 else
"111111110000" when X = 9 AND Y = 28 else
"111111110000" when X = 10 AND Y = 28 else
"111111110000" when X = 11 AND Y = 28 else
"111111110000" when X = 12 AND Y = 28 else
"111111110000" when X = 13 AND Y = 28 else
"111111110000" when X = 14 AND Y = 28 else
"111111110000" when X = 15 AND Y = 28 else
"111111110000" when X = 16 AND Y = 28 else
"111111110000" when X = 17 AND Y = 28 else
"111111110000" when X = 18 AND Y = 28 else
"111111110000" when X = 19 AND Y = 28 else
"111111110000" when X = 20 AND Y = 28 else
"111111110000" when X = 21 AND Y = 28 else
"111111110000" when X = 22 AND Y = 28 else
"111111110000" when X = 23 AND Y = 28 else
"111111110000" when X = 24 AND Y = 28 else
"111111110000" when X = 25 AND Y = 28 else
"111111110000" when X = 26 AND Y = 28 else
"111111110000" when X = 27 AND Y = 28 else
"111111110000" when X = 28 AND Y = 28 else
"111111110000" when X = 29 AND Y = 28 else
"111111110000" when X = 30 AND Y = 28 else
"111111110000" when X = 31 AND Y = 28 else
"111111110000" when X = 32 AND Y = 28 else
"111111110000" when X = 33 AND Y = 28 else
"111111110000" when X = 34 AND Y = 28 else
"111111110000" when X = 35 AND Y = 28 else
"111111110000" when X = 36 AND Y = 28 else
"111111110000" when X = 37 AND Y = 28 else
"111111110000" when X = 38 AND Y = 28 else
"111111110000" when X = 39 AND Y = 28 else
"111111110000" when X = 40 AND Y = 28 else
"111111110000" when X = 41 AND Y = 28 else
"111111110000" when X = 42 AND Y = 28 else
"111111110000" when X = 43 AND Y = 28 else
"111111110000" when X = 44 AND Y = 28 else
"111111110000" when X = 45 AND Y = 28 else
"111111110000" when X = 0 AND Y = 29 else
"111111110000" when X = 1 AND Y = 29 else
"111111110000" when X = 2 AND Y = 29 else
"111111110000" when X = 3 AND Y = 29 else
"111111110000" when X = 4 AND Y = 29 else
"111111110000" when X = 5 AND Y = 29 else
"111111110000" when X = 6 AND Y = 29 else
"111111110000" when X = 7 AND Y = 29 else
"111111110000" when X = 8 AND Y = 29 else
"111111110000" when X = 9 AND Y = 29 else
"111111110000" when X = 10 AND Y = 29 else
"111111110000" when X = 11 AND Y = 29 else
"111111110000" when X = 12 AND Y = 29 else
"111111110000" when X = 13 AND Y = 29 else
"111111110000" when X = 14 AND Y = 29 else
"111111110000" when X = 15 AND Y = 29 else
"111111110000" when X = 16 AND Y = 29 else
"111111110000" when X = 17 AND Y = 29 else
"111111110000" when X = 18 AND Y = 29 else
"111111110000" when X = 19 AND Y = 29 else
"111111110000" when X = 20 AND Y = 29 else
"111111110000" when X = 21 AND Y = 29 else
"111111110000" when X = 22 AND Y = 29 else
"111111110000" when X = 23 AND Y = 29 else
"111111110000" when X = 24 AND Y = 29 else
"111111110000" when X = 25 AND Y = 29 else
"111111110000" when X = 26 AND Y = 29 else
"111111110000" when X = 27 AND Y = 29 else
"111111110000" when X = 28 AND Y = 29 else
"111111110000" when X = 29 AND Y = 29 else
"111111110000" when X = 30 AND Y = 29 else
"111111110000" when X = 31 AND Y = 29 else
"111111110000" when X = 32 AND Y = 29 else
"111111110000" when X = 33 AND Y = 29 else
"111111110000" when X = 34 AND Y = 29 else
"111111110000" when X = 35 AND Y = 29 else
"111111110000" when X = 36 AND Y = 29 else
"111111110000" when X = 37 AND Y = 29 else
"111111110000" when X = 38 AND Y = 29 else
"111111110000" when X = 39 AND Y = 29 else
"111111110000" when X = 40 AND Y = 29 else
"111111110000" when X = 41 AND Y = 29 else
"111111110000" when X = 42 AND Y = 29 else
"111111110000" when X = 43 AND Y = 29 else
"111111110000" when X = 44 AND Y = 29 else
"111111110000" when X = 45 AND Y = 29 else
"000000000000"; -- should never get here
end rtl;
