-- Tyler Hansen
-- CS232 Final Project
-- genSpriteROM.py
-- generates a ROM file in VHDL from a .ppm image

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity player_sprite is
port(
X	: in INTEGER RANGE 0 TO 1688;
Y	: in INTEGER RANGE 0 TO 1688;
data : out std_logic_vector (11 downto 0)
);

end entity;

architecture rtl of player_sprite is
begin
data <=
"111111110000" when X = 0 AND Y = 0 else "111111110000" when X = 1 AND Y = 0 else "111111110000" when X = 2 AND Y = 0 else "111111110000" when X = 3 AND Y = 0 else "111111110000" when X = 4 AND Y = 0 else "111111110000" when X = 5 AND Y = 0 else "111111110000" when X = 6 AND Y = 0 else "111111110000" when X = 7 AND Y = 0 else "111111110000" when X = 8 AND Y = 0 else "111111110000" when X = 9 AND Y = 0 else "111111110000" when X = 10 AND Y = 0 else "111111110000" when X = 11 AND Y = 0 else "111111110000" when X = 12 AND Y = 0 else "111111110000" when X = 13 AND Y = 0 else "111111110000" when X = 14 AND Y = 0 else "111111110000" when X = 15 AND Y = 0 else "111111110000" when X = 16 AND Y = 0 else "111111110000" when X = 17 AND Y = 0 else "111111110000" when X = 18 AND Y = 0 else "111111110000" when X = 19 AND Y = 0 else "111111110000" when X = 20 AND Y = 0 else "111111110000" when X = 21 AND Y = 0 else "111111110000" when X = 22 AND Y = 0 else "111111110000" when X = 23 AND Y = 0 else "111111110000" when X = 24 AND Y = 0 else "111111110000" when X = 25 AND Y = 0 else "111111110000" when X = 26 AND Y = 0 else "111111110000" when X = 27 AND Y = 0 else "111111110000" when X = 28 AND Y = 0 else "111111110000" when X = 29 AND Y = 0 else "111111110000" when X = 30 AND Y = 0 else "111111110000" when X = 31 AND Y = 0 else "111111110000" when X = 32 AND Y = 0 else "111111110000" when X = 33 AND Y = 0 else "111111110000" when X = 34 AND Y = 0 else "111111110000" when X = 35 AND Y = 0 else "111111110000" when X = 36 AND Y = 0 else "111111110000" when X = 37 AND Y = 0 else "111111110000" when X = 38 AND Y = 0 else "111111110000" when X = 39 AND Y = 0 else "111111110000" when X = 40 AND Y = 0 else "111111110000" when X = 41 AND Y = 0 else "111111110000" when X = 42 AND Y = 0 else "111111110000" when X = 43 AND Y = 0 else "111111110000" when X = 44 AND Y = 0 else "111111110000" when X = 45 AND Y = 0 else "111111110000" when X = 46 AND Y = 0 else "111111110000" when X = 47 AND Y = 0 else "111111110000" when X = 48 AND Y = 0 else "111111110000" when X = 49 AND Y = 0 else "111111110000" when X = 50 AND Y = 0 else "111111110000" when X = 51 AND Y = 0 else "111111110000" when X = 52 AND Y = 0 else "111111110000" when X = 53 AND Y = 0 else "111111110000" when X = 54 AND Y = 0 else "111111110000" when X = 55 AND Y = 0 else "111111110000" when X = 56 AND Y = 0 else "111111110000" when X = 57 AND Y = 0 else "111111110000" when X = 58 AND Y = 0 else "111111110000" when X = 59 AND Y = 0 else "111111110000" when X = 60 AND Y = 0 else "111111110000" when X = 61 AND Y = 0 else "111111110000" when X = 62 AND Y = 0 else "111111110000" when X = 63 AND Y = 0 else "111111110000" when X = 64 AND Y = 0 else "111111110000" when X = 65 AND Y = 0 else "111111110000" when X = 66 AND Y = 0 else "111111110000" when X = 67 AND Y = 0 else "111111110000" when X = 68 AND Y = 0 else "111111110000" when X = 0 AND Y = 1 else "111111110000" when X = 1 AND Y = 1 else "111111110000" when X = 2 AND Y = 1 else "111111110000" when X = 3 AND Y = 1 else "111111110000" when X = 4 AND Y = 1 else "111111110000" when X = 5 AND Y = 1 else "111111110000" when X = 6 AND Y = 1 else "111111110000" when X = 7 AND Y = 1 else "111111110000" when X = 8 AND Y = 1 else "111111110000" when X = 9 AND Y = 1 else "111111110000" when X = 10 AND Y = 1 else "111111110000" when X = 11 AND Y = 1 else "111111110000" when X = 12 AND Y = 1 else "111111110000" when X = 13 AND Y = 1 else "111111110000" when X = 14 AND Y = 1 else "111111110000" when X = 15 AND Y = 1 else "111111110000" when X = 16 AND Y = 1 else "111111110000" when X = 17 AND Y = 1 else "111111110000" when X = 18 AND Y = 1 else "111111110000" when X = 19 AND Y = 1 else "111111110000" when X = 20 AND Y = 1 else "111111110000" when X = 21 AND Y = 1 else "111111110000" when X = 22 AND Y = 1 else "111111110000" when X = 23 AND Y = 1 else "111111110000" when X = 24 AND Y = 1 else "111111110000" when X = 25 AND Y = 1 else "111111110000" when X = 26 AND Y = 1 else "111111110000" when X = 27 AND Y = 1 else "111111110000" when X = 28 AND Y = 1 else "111111110000" when X = 29 AND Y = 1 else "111111110000" when X = 30 AND Y = 1 else "111111110000" when X = 31 AND Y = 1 else "111111110000" when X = 32 AND Y = 1 else "111111110000" when X = 33 AND Y = 1 else "111111110000" when X = 34 AND Y = 1 else "111111110000" when X = 35 AND Y = 1 else "111111110000" when X = 36 AND Y = 1 else "111111110000" when X = 37 AND Y = 1 else "111111110000" when X = 38 AND Y = 1 else "111111110000" when X = 39 AND Y = 1 else "111111110000" when X = 40 AND Y = 1 else "111111110000" when X = 41 AND Y = 1 else "111111110000" when X = 42 AND Y = 1 else "111111110000" when X = 43 AND Y = 1 else "111111110000" when X = 44 AND Y = 1 else "111111110000" when X = 45 AND Y = 1 else "111111110000" when X = 46 AND Y = 1 else "111111110000" when X = 47 AND Y = 1 else "111111110000" when X = 48 AND Y = 1 else "111111110000" when X = 49 AND Y = 1 else "111111110000" when X = 50 AND Y = 1 else "111111110000" when X = 51 AND Y = 1 else "111111110000" when X = 52 AND Y = 1 else "111111110000" when X = 53 AND Y = 1 else "111111110000" when X = 54 AND Y = 1 else "111111110000" when X = 55 AND Y = 1 else "111111110000" when X = 56 AND Y = 1 else "111111110000" when X = 57 AND Y = 1 else "111111110000" when X = 58 AND Y = 1 else "111111110000" when X = 59 AND Y = 1 else "111111110000" when X = 60 AND Y = 1 else "111111110000" when X = 61 AND Y = 1 else "111111110000" when X = 62 AND Y = 1 else "111111110000" when X = 63 AND Y = 1 else "111111110000" when X = 64 AND Y = 1 else "111111110000" when X = 65 AND Y = 1 else "111111110000" when X = 66 AND Y = 1 else "111111110000" when X = 67 AND Y = 1 else "111111110000" when X = 68 AND Y = 1 else "111111110000" when X = 0 AND Y = 2 else "111111110000" when X = 1 AND Y = 2 else "111111110000" when X = 2 AND Y = 2 else "111111110000" when X = 3 AND Y = 2 else "111111110000" when X = 4 AND Y = 2 else "111111110000" when X = 5 AND Y = 2 else "111111110000" when X = 6 AND Y = 2 else "111111110000" when X = 7 AND Y = 2 else "111111110000" when X = 8 AND Y = 2 else "111111110000" when X = 9 AND Y = 2 else "111111110000" when X = 10 AND Y = 2 else "111111110000" when X = 11 AND Y = 2 else "111111110000" when X = 12 AND Y = 2 else "111111110000" when X = 13 AND Y = 2 else "111111110000" when X = 14 AND Y = 2 else "111111110000" when X = 15 AND Y = 2 else "111111110000" when X = 16 AND Y = 2 else "111111110000" when X = 17 AND Y = 2 else "111111110000" when X = 18 AND Y = 2 else "111111110000" when X = 19 AND Y = 2 else "111111110000" when X = 20 AND Y = 2 else "111111110000" when X = 21 AND Y = 2 else "111111110000" when X = 22 AND Y = 2 else "111111110000" when X = 23 AND Y = 2 else "111111110000" when X = 24 AND Y = 2 else "111111110000" when X = 25 AND Y = 2 else "111111110000" when X = 26 AND Y = 2 else "111111110000" when X = 27 AND Y = 2 else "111111110000" when X = 28 AND Y = 2 else "111111110000" when X = 29 AND Y = 2 else "111111110000" when X = 30 AND Y = 2 else "111111110000" when X = 31 AND Y = 2 else "111111110000" when X = 32 AND Y = 2 else "111111110000" when X = 33 AND Y = 2 else "111111110000" when X = 34 AND Y = 2 else "111111110000" when X = 35 AND Y = 2 else "111111110000" when X = 36 AND Y = 2 else "111111110000" when X = 37 AND Y = 2 else "111111110000" when X = 38 AND Y = 2 else "111111110000" when X = 39 AND Y = 2 else "111111110000" when X = 40 AND Y = 2 else "111111110000" when X = 41 AND Y = 2 else "111111110000" when X = 42 AND Y = 2 else "111111110000" when X = 43 AND Y = 2 else "111111110000" when X = 44 AND Y = 2 else "111111110000" when X = 45 AND Y = 2 else "111111110000" when X = 46 AND Y = 2 else "111111110000" when X = 47 AND Y = 2 else "111111110000" when X = 48 AND Y = 2 else "111111110000" when X = 49 AND Y = 2 else "111111110000" when X = 50 AND Y = 2 else "111111110000" when X = 51 AND Y = 2 else "111111110000" when X = 52 AND Y = 2 else "111111110000" when X = 53 AND Y = 2 else "111111110000" when X = 54 AND Y = 2 else "111111110000" when X = 55 AND Y = 2 else "111111110000" when X = 56 AND Y = 2 else "111111110000" when X = 57 AND Y = 2 else "111111110000" when X = 58 AND Y = 2 else "111111110000" when X = 59 AND Y = 2 else "111111110000" when X = 60 AND Y = 2 else "111111110000" when X = 61 AND Y = 2 else "111111110000" when X = 62 AND Y = 2 else "111111110000" when X = 63 AND Y = 2 else "111111110000" when X = 64 AND Y = 2 else "111111110000" when X = 65 AND Y = 2 else "111111110000" when X = 66 AND Y = 2 else "111111110000" when X = 67 AND Y = 2 else "111111110000" when X = 68 AND Y = 2 else "111111110000" when X = 0 AND Y = 3 else "111111110000" when X = 1 AND Y = 3 else "111111110000" when X = 2 AND Y = 3 else "111111110000" when X = 3 AND Y = 3 else "111111110000" when X = 4 AND Y = 3 else "111111110000" when X = 5 AND Y = 3 else "111111110000" when X = 6 AND Y = 3 else "111111110000" when X = 7 AND Y = 3 else "111111110000" when X = 8 AND Y = 3 else "111111110000" when X = 9 AND Y = 3 else "111111110000" when X = 10 AND Y = 3 else "111111110000" when X = 11 AND Y = 3 else "111111110000" when X = 12 AND Y = 3 else "111111110000" when X = 13 AND Y = 3 else "111111110000" when X = 14 AND Y = 3 else "111111110000" when X = 15 AND Y = 3 else "111111110000" when X = 16 AND Y = 3 else "111111110000" when X = 17 AND Y = 3 else "111111110000" when X = 18 AND Y = 3 else "111111110000" when X = 19 AND Y = 3 else "111111110000" when X = 20 AND Y = 3 else "111111110000" when X = 21 AND Y = 3 else "111111110000" when X = 22 AND Y = 3 else "111111110000" when X = 23 AND Y = 3 else "111111110000" when X = 24 AND Y = 3 else "111111110000" when X = 25 AND Y = 3 else "111111110000" when X = 26 AND Y = 3 else "111111110000" when X = 27 AND Y = 3 else "111111110000" when X = 28 AND Y = 3 else "111111110000" when X = 29 AND Y = 3 else "111111110000" when X = 30 AND Y = 3 else "111111110000" when X = 31 AND Y = 3 else "111111110000" when X = 32 AND Y = 3 else "111111110000" when X = 33 AND Y = 3 else "111111110000" when X = 34 AND Y = 3 else "111111110000" when X = 35 AND Y = 3 else "111111110000" when X = 36 AND Y = 3 else "111111110000" when X = 37 AND Y = 3 else "111111110000" when X = 38 AND Y = 3 else "111111110000" when X = 39 AND Y = 3 else "111111110000" when X = 40 AND Y = 3 else "111111110000" when X = 41 AND Y = 3 else "111111110000" when X = 42 AND Y = 3 else "111111110000" when X = 43 AND Y = 3 else "111111110000" when X = 44 AND Y = 3 else "111111110000" when X = 45 AND Y = 3 else "111111110000" when X = 46 AND Y = 3 else "111111110000" when X = 47 AND Y = 3 else "111111110000" when X = 48 AND Y = 3 else "111111110000" when X = 49 AND Y = 3 else "111111110000" when X = 50 AND Y = 3 else "111111110000" when X = 51 AND Y = 3 else "111111110000" when X = 52 AND Y = 3 else "111111110000" when X = 53 AND Y = 3 else "111111110000" when X = 54 AND Y = 3 else "111111110000" when X = 55 AND Y = 3 else "111111110000" when X = 56 AND Y = 3 else "111111110000" when X = 57 AND Y = 3 else "111111110000" when X = 58 AND Y = 3 else "111111110000" when X = 59 AND Y = 3 else "111111110000" when X = 60 AND Y = 3 else "111111110000" when X = 61 AND Y = 3 else "111111110000" when X = 62 AND Y = 3 else "111111110000" when X = 63 AND Y = 3 else "111111110000" when X = 64 AND Y = 3 else "111111110000" when X = 65 AND Y = 3 else "111111110000" when X = 66 AND Y = 3 else "111111110000" when X = 67 AND Y = 3 else "111111110000" when X = 68 AND Y = 3 else "111111110000" when X = 0 AND Y = 4 else "111111110000" when X = 1 AND Y = 4 else "111111110000" when X = 2 AND Y = 4 else "111111110000" when X = 3 AND Y = 4 else "111111110000" when X = 4 AND Y = 4 else "111111110000" when X = 5 AND Y = 4 else "111111110000" when X = 6 AND Y = 4 else "111111110000" when X = 7 AND Y = 4 else "111111110000" when X = 8 AND Y = 4 else "111111110000" when X = 9 AND Y = 4 else "111111110000" when X = 10 AND Y = 4 else "111111110000" when X = 11 AND Y = 4 else "111111110000" when X = 12 AND Y = 4 else "111111110000" when X = 13 AND Y = 4 else "111111110000" when X = 14 AND Y = 4 else "111111110000" when X = 15 AND Y = 4 else "111111110000" when X = 16 AND Y = 4 else "111111110000" when X = 17 AND Y = 4 else "111111110000" when X = 18 AND Y = 4 else "111111110000" when X = 19 AND Y = 4 else "111111110000" when X = 20 AND Y = 4 else "111111110000" when X = 21 AND Y = 4 else "111111110000" when X = 22 AND Y = 4 else "111111110000" when X = 23 AND Y = 4 else "111111110000" when X = 24 AND Y = 4 else "111111110000" when X = 25 AND Y = 4 else "111111110000" when X = 26 AND Y = 4 else "111111110000" when X = 27 AND Y = 4 else "111111110000" when X = 28 AND Y = 4 else "111111110000" when X = 29 AND Y = 4 else "111111110000" when X = 30 AND Y = 4 else "111111110000" when X = 31 AND Y = 4 else "111111110101" when X = 32 AND Y = 4 else "111111110101" when X = 33 AND Y = 4 else "111111110101" when X = 34 AND Y = 4 else "111111110000" when X = 35 AND Y = 4 else "111111110000" when X = 36 AND Y = 4 else "111111110000" when X = 37 AND Y = 4 else "111111110000" when X = 38 AND Y = 4 else "111111110000" when X = 39 AND Y = 4 else "111111110000" when X = 40 AND Y = 4 else "111111110000" when X = 41 AND Y = 4 else "111111110000" when X = 42 AND Y = 4 else "111111110000" when X = 43 AND Y = 4 else "111111110000" when X = 44 AND Y = 4 else "111111110000" when X = 45 AND Y = 4 else "111111110000" when X = 46 AND Y = 4 else "111111110000" when X = 47 AND Y = 4 else "111111110000" when X = 48 AND Y = 4 else "111111110000" when X = 49 AND Y = 4 else "111111110000" when X = 50 AND Y = 4 else "111111110000" when X = 51 AND Y = 4 else "111111110000" when X = 52 AND Y = 4 else "111111110000" when X = 53 AND Y = 4 else "111111110000" when X = 54 AND Y = 4 else "111111110000" when X = 55 AND Y = 4 else "111111110000" when X = 56 AND Y = 4 else "111111110000" when X = 57 AND Y = 4 else "111111110000" when X = 58 AND Y = 4 else "111111110000" when X = 59 AND Y = 4 else "111111110000" when X = 60 AND Y = 4 else "111111110000" when X = 61 AND Y = 4 else "111111110000" when X = 62 AND Y = 4 else "111111110000" when X = 63 AND Y = 4 else "111111110000" when X = 64 AND Y = 4 else "111111110000" when X = 65 AND Y = 4 else "111111110000" when X = 66 AND Y = 4 else "111111110000" when X = 67 AND Y = 4 else "111111110000" when X = 68 AND Y = 4 else "111111110000" when X = 0 AND Y = 5 else "111111110000" when X = 1 AND Y = 5 else "111111110000" when X = 2 AND Y = 5 else "111111110000" when X = 3 AND Y = 5 else "111111110000" when X = 4 AND Y = 5 else "111111110000" when X = 5 AND Y = 5 else "111111110000" when X = 6 AND Y = 5 else "111111110000" when X = 7 AND Y = 5 else "111111110000" when X = 8 AND Y = 5 else "111111110000" when X = 9 AND Y = 5 else "111111110000" when X = 10 AND Y = 5 else "111111110000" when X = 11 AND Y = 5 else "111111110000" when X = 12 AND Y = 5 else "111111110000" when X = 13 AND Y = 5 else "111111110000" when X = 14 AND Y = 5 else "111111110000" when X = 15 AND Y = 5 else "111111110000" when X = 16 AND Y = 5 else "111111110000" when X = 17 AND Y = 5 else "111111110000" when X = 18 AND Y = 5 else "111111110000" when X = 19 AND Y = 5 else "111111110000" when X = 20 AND Y = 5 else "111111110000" when X = 21 AND Y = 5 else "111111110000" when X = 22 AND Y = 5 else "111111110000" when X = 23 AND Y = 5 else "111111110000" when X = 24 AND Y = 5 else "111111110000" when X = 25 AND Y = 5 else "111111110000" when X = 26 AND Y = 5 else "111111110000" when X = 27 AND Y = 5 else "111111110000" when X = 28 AND Y = 5 else "111111110000" when X = 29 AND Y = 5 else "111111110000" when X = 30 AND Y = 5 else "001101101111" when X = 31 AND Y = 5 else "000100111111" when X = 32 AND Y = 5 else "000100111111" when X = 33 AND Y = 5 else "000100111111" when X = 34 AND Y = 5 else "001001001111" when X = 35 AND Y = 5 else "101011011101" when X = 36 AND Y = 5 else "111111110000" when X = 37 AND Y = 5 else "111111110000" when X = 38 AND Y = 5 else "111111110000" when X = 39 AND Y = 5 else "111111110000" when X = 40 AND Y = 5 else "111111110000" when X = 41 AND Y = 5 else "111111110000" when X = 42 AND Y = 5 else "111111110000" when X = 43 AND Y = 5 else "111111110000" when X = 44 AND Y = 5 else "111111110000" when X = 45 AND Y = 5 else "111111110000" when X = 46 AND Y = 5 else "111111110000" when X = 47 AND Y = 5 else "111111110000" when X = 48 AND Y = 5 else "111111110000" when X = 49 AND Y = 5 else "111111110000" when X = 50 AND Y = 5 else "111111110000" when X = 51 AND Y = 5 else "111111110000" when X = 52 AND Y = 5 else "111111110000" when X = 53 AND Y = 5 else "111111110000" when X = 54 AND Y = 5 else "111111110000" when X = 55 AND Y = 5 else "111111110000" when X = 56 AND Y = 5 else "111111110000" when X = 57 AND Y = 5 else "111111110000" when X = 58 AND Y = 5 else "111111110000" when X = 59 AND Y = 5 else "111111110000" when X = 60 AND Y = 5 else "111111110000" when X = 61 AND Y = 5 else "111111110000" when X = 62 AND Y = 5 else "111111110000" when X = 63 AND Y = 5 else "111111110000" when X = 64 AND Y = 5 else "111111110000" when X = 65 AND Y = 5 else "111111110000" when X = 66 AND Y = 5 else "111111110000" when X = 67 AND Y = 5 else "111111110000" when X = 68 AND Y = 5 else "111111110000" when X = 0 AND Y = 6 else "111111110000" when X = 1 AND Y = 6 else "111111110000" when X = 2 AND Y = 6 else "111111110000" when X = 3 AND Y = 6 else "111111110000" when X = 4 AND Y = 6 else "111111110000" when X = 5 AND Y = 6 else "111111110000" when X = 6 AND Y = 6 else "111111110000" when X = 7 AND Y = 6 else "111111110000" when X = 8 AND Y = 6 else "111111110000" when X = 9 AND Y = 6 else "111111110000" when X = 10 AND Y = 6 else "111111110000" when X = 11 AND Y = 6 else "111111110000" when X = 12 AND Y = 6 else "111111110000" when X = 13 AND Y = 6 else "111111110000" when X = 14 AND Y = 6 else "111111110000" when X = 15 AND Y = 6 else "111111110000" when X = 16 AND Y = 6 else "111111110000" when X = 17 AND Y = 6 else "111111110000" when X = 18 AND Y = 6 else "111111110000" when X = 19 AND Y = 6 else "111111110000" when X = 20 AND Y = 6 else "111111110000" when X = 21 AND Y = 6 else "111111110000" when X = 22 AND Y = 6 else "111111110000" when X = 23 AND Y = 6 else "111111110000" when X = 24 AND Y = 6 else "111111110000" when X = 25 AND Y = 6 else "111111110000" when X = 26 AND Y = 6 else "111111110000" when X = 27 AND Y = 6 else "111111110000" when X = 28 AND Y = 6 else "111111110000" when X = 29 AND Y = 6 else "001101101111" when X = 30 AND Y = 6 else "000100011111" when X = 31 AND Y = 6 else "001101101111" when X = 32 AND Y = 6 else "011010011111" when X = 33 AND Y = 6 else "010001111111" when X = 34 AND Y = 6 else "000100011111" when X = 35 AND Y = 6 else "001001011111" when X = 36 AND Y = 6 else "100010111110" when X = 37 AND Y = 6 else "111111110000" when X = 38 AND Y = 6 else "111111110000" when X = 39 AND Y = 6 else "111111110000" when X = 40 AND Y = 6 else "111111110000" when X = 41 AND Y = 6 else "111111110000" when X = 42 AND Y = 6 else "111111110000" when X = 43 AND Y = 6 else "111111110000" when X = 44 AND Y = 6 else "111111110000" when X = 45 AND Y = 6 else "111111110000" when X = 46 AND Y = 6 else "111111110000" when X = 47 AND Y = 6 else "111111110000" when X = 48 AND Y = 6 else "111111110000" when X = 49 AND Y = 6 else "111111110000" when X = 50 AND Y = 6 else "111111110000" when X = 51 AND Y = 6 else "111111110000" when X = 52 AND Y = 6 else "111111110000" when X = 53 AND Y = 6 else "111111110000" when X = 54 AND Y = 6 else "111111110000" when X = 55 AND Y = 6 else "111111110000" when X = 56 AND Y = 6 else "111111110000" when X = 57 AND Y = 6 else "111111110000" when X = 58 AND Y = 6 else "111111110000" when X = 59 AND Y = 6 else "111111110000" when X = 60 AND Y = 6 else "111111110000" when X = 61 AND Y = 6 else "111111110000" when X = 62 AND Y = 6 else "111111110000" when X = 63 AND Y = 6 else "111111110000" when X = 64 AND Y = 6 else "111111110000" when X = 65 AND Y = 6 else "111111110000" when X = 66 AND Y = 6 else "111111110000" when X = 67 AND Y = 6 else "111111110000" when X = 68 AND Y = 6 else "111111110000" when X = 0 AND Y = 7 else "111111110000" when X = 1 AND Y = 7 else "111111110000" when X = 2 AND Y = 7 else "111111110000" when X = 3 AND Y = 7 else "111111110000" when X = 4 AND Y = 7 else "111111110000" when X = 5 AND Y = 7 else "111111110000" when X = 6 AND Y = 7 else "111111110000" when X = 7 AND Y = 7 else "111111110000" when X = 8 AND Y = 7 else "111111110000" when X = 9 AND Y = 7 else "111111110000" when X = 10 AND Y = 7 else "111111110000" when X = 11 AND Y = 7 else "111111110000" when X = 12 AND Y = 7 else "111111110000" when X = 13 AND Y = 7 else "111111110000" when X = 14 AND Y = 7 else "111111110000" when X = 15 AND Y = 7 else "111111110000" when X = 16 AND Y = 7 else "111111110000" when X = 17 AND Y = 7 else "111111110000" when X = 18 AND Y = 7 else "111111110000" when X = 19 AND Y = 7 else "111111110000" when X = 20 AND Y = 7 else "111111110000" when X = 21 AND Y = 7 else "111111110000" when X = 22 AND Y = 7 else "111111110000" when X = 23 AND Y = 7 else "111111110000" when X = 24 AND Y = 7 else "111111110000" when X = 25 AND Y = 7 else "111111110000" when X = 26 AND Y = 7 else "111111110000" when X = 27 AND Y = 7 else "100111001110" when X = 28 AND Y = 7 else "010001111111" when X = 29 AND Y = 7 else "000100011111" when X = 30 AND Y = 7 else "000001011111" when X = 31 AND Y = 7 else "001110111110" when X = 32 AND Y = 7 else "011011011110" when X = 33 AND Y = 7 else "010011001110" when X = 34 AND Y = 7 else "000001101110" when X = 35 AND Y = 7 else "000100011111" when X = 36 AND Y = 7 else "001101101111" when X = 37 AND Y = 7 else "011110111111" when X = 38 AND Y = 7 else "111111110000" when X = 39 AND Y = 7 else "111111110000" when X = 40 AND Y = 7 else "111111110000" when X = 41 AND Y = 7 else "111111110000" when X = 42 AND Y = 7 else "111111110000" when X = 43 AND Y = 7 else "111111110000" when X = 44 AND Y = 7 else "111111110000" when X = 45 AND Y = 7 else "111111110000" when X = 46 AND Y = 7 else "111111110000" when X = 47 AND Y = 7 else "111111110000" when X = 48 AND Y = 7 else "111111110000" when X = 49 AND Y = 7 else "111111110000" when X = 50 AND Y = 7 else "111111110000" when X = 51 AND Y = 7 else "111111110000" when X = 52 AND Y = 7 else "111111110000" when X = 53 AND Y = 7 else "111111110000" when X = 54 AND Y = 7 else "111111110000" when X = 55 AND Y = 7 else "111111110000" when X = 56 AND Y = 7 else "111111110000" when X = 57 AND Y = 7 else "111111110000" when X = 58 AND Y = 7 else "111111110000" when X = 59 AND Y = 7 else "111111110000" when X = 60 AND Y = 7 else "111111110000" when X = 61 AND Y = 7 else "111111110000" when X = 62 AND Y = 7 else "111111110000" when X = 63 AND Y = 7 else "111111110000" when X = 64 AND Y = 7 else "111111110000" when X = 65 AND Y = 7 else "111111110000" when X = 66 AND Y = 7 else "111111110000" when X = 67 AND Y = 7 else "111111110000" when X = 68 AND Y = 7 else "111111110000" when X = 0 AND Y = 8 else "111111110000" when X = 1 AND Y = 8 else "111111110000" when X = 2 AND Y = 8 else "111111110000" when X = 3 AND Y = 8 else "111111110000" when X = 4 AND Y = 8 else "111111110000" when X = 5 AND Y = 8 else "111111110000" when X = 6 AND Y = 8 else "111111110000" when X = 7 AND Y = 8 else "111111110000" when X = 8 AND Y = 8 else "111111110000" when X = 9 AND Y = 8 else "100011001101" when X = 10 AND Y = 8 else "011010011001" when X = 11 AND Y = 8 else "011010011001" when X = 12 AND Y = 8 else "011010011001" when X = 13 AND Y = 8 else "011010011001" when X = 14 AND Y = 8 else "011110101011" when X = 15 AND Y = 8 else "111111110000" when X = 16 AND Y = 8 else "111111110000" when X = 17 AND Y = 8 else "111111110000" when X = 18 AND Y = 8 else "111111110000" when X = 19 AND Y = 8 else "111111110000" when X = 20 AND Y = 8 else "111111110000" when X = 21 AND Y = 8 else "111111110000" when X = 22 AND Y = 8 else "111111110000" when X = 23 AND Y = 8 else "101111001011" when X = 24 AND Y = 8 else "101111001010" when X = 25 AND Y = 8 else "110010111010" when X = 26 AND Y = 8 else "101010111011" when X = 27 AND Y = 8 else "010110111110" when X = 28 AND Y = 8 else "000100011111" when X = 29 AND Y = 8 else "000100001111" when X = 30 AND Y = 8 else "010110101011" when X = 31 AND Y = 8 else "011111101001" when X = 32 AND Y = 8 else "011111011010" when X = 33 AND Y = 8 else "011111011010" when X = 34 AND Y = 8 else "011011001010" when X = 35 AND Y = 8 else "000100101111" when X = 36 AND Y = 8 else "000100001111" when X = 37 AND Y = 8 else "010010001111" when X = 38 AND Y = 8 else "100111001100" when X = 39 AND Y = 8 else "110010101010" when X = 40 AND Y = 8 else "101110111010" when X = 41 AND Y = 8 else "101111001010" when X = 42 AND Y = 8 else "101011011101" when X = 43 AND Y = 8 else "111111110000" when X = 44 AND Y = 8 else "111111110000" when X = 45 AND Y = 8 else "111111110000" when X = 46 AND Y = 8 else "111111110000" when X = 47 AND Y = 8 else "111111110000" when X = 48 AND Y = 8 else "111111110000" when X = 49 AND Y = 8 else "111111110000" when X = 50 AND Y = 8 else "100011001101" when X = 51 AND Y = 8 else "011010011010" when X = 52 AND Y = 8 else "011010011001" when X = 53 AND Y = 8 else "011010011001" when X = 54 AND Y = 8 else "011010011001" when X = 55 AND Y = 8 else "100010111100" when X = 56 AND Y = 8 else "111111110000" when X = 57 AND Y = 8 else "111111110000" when X = 58 AND Y = 8 else "111111110000" when X = 59 AND Y = 8 else "111111110000" when X = 60 AND Y = 8 else "111111110000" when X = 61 AND Y = 8 else "111111110000" when X = 62 AND Y = 8 else "111111110000" when X = 63 AND Y = 8 else "111111110000" when X = 64 AND Y = 8 else "111111110000" when X = 65 AND Y = 8 else "111111110000" when X = 66 AND Y = 8 else "111111110000" when X = 67 AND Y = 8 else "111111110000" when X = 68 AND Y = 8 else "111111110000" when X = 0 AND Y = 9 else "111111110000" when X = 1 AND Y = 9 else "111111110000" when X = 2 AND Y = 9 else "111111110000" when X = 3 AND Y = 9 else "111111110000" when X = 4 AND Y = 9 else "111111110000" when X = 5 AND Y = 9 else "111111110000" when X = 6 AND Y = 9 else "111111110000" when X = 7 AND Y = 9 else "111111110000" when X = 8 AND Y = 9 else "101011011100" when X = 9 AND Y = 9 else "010110001000" when X = 10 AND Y = 9 else "000100010001" when X = 11 AND Y = 9 else "000100010001" when X = 12 AND Y = 9 else "000000000000" when X = 13 AND Y = 9 else "000000000000" when X = 14 AND Y = 9 else "001000110011" when X = 15 AND Y = 9 else "011110111100" when X = 16 AND Y = 9 else "111111110000" when X = 17 AND Y = 9 else "111111110000" when X = 18 AND Y = 9 else "100111001110" when X = 19 AND Y = 9 else "100110111101" when X = 20 AND Y = 9 else "100110111101" when X = 21 AND Y = 9 else "100110111101" when X = 22 AND Y = 9 else "101111001011" when X = 23 AND Y = 9 else "111110010011" when X = 24 AND Y = 9 else "111110000000" when X = 25 AND Y = 9 else "111101000000" when X = 26 AND Y = 9 else "110001100101" when X = 27 AND Y = 9 else "000010101101" when X = 28 AND Y = 9 else "000100011111" when X = 29 AND Y = 9 else "000100001111" when X = 30 AND Y = 9 else "101010110111" when X = 31 AND Y = 9 else "111111110000" when X = 32 AND Y = 9 else "111111110000" when X = 33 AND Y = 9 else "111111110000" when X = 34 AND Y = 9 else "110111010100" when X = 35 AND Y = 9 else "000100101110" when X = 36 AND Y = 9 else "000100001111" when X = 37 AND Y = 9 else "000010011110" when X = 38 AND Y = 9 else "101010001000" when X = 39 AND Y = 9 else "111100010000" when X = 40 AND Y = 9 else "111101110000" when X = 41 AND Y = 9 else "111110000000" when X = 42 AND Y = 9 else "110110111000" when X = 43 AND Y = 9 else "101011001101" when X = 44 AND Y = 9 else "100110111101" when X = 45 AND Y = 9 else "100110111101" when X = 46 AND Y = 9 else "100110111101" when X = 47 AND Y = 9 else "111111110000" when X = 48 AND Y = 9 else "111111110000" when X = 49 AND Y = 9 else "110011101010" when X = 50 AND Y = 9 else "010110001000" when X = 51 AND Y = 9 else "000000000000" when X = 52 AND Y = 9 else "000000000000" when X = 53 AND Y = 9 else "000100010001" when X = 54 AND Y = 9 else "000100010001" when X = 55 AND Y = 9 else "010001100110" when X = 56 AND Y = 9 else "100011001101" when X = 57 AND Y = 9 else "111111110000" when X = 58 AND Y = 9 else "111111110000" when X = 59 AND Y = 9 else "111111110000" when X = 60 AND Y = 9 else "111111110000" when X = 61 AND Y = 9 else "111111110000" when X = 62 AND Y = 9 else "111111110000" when X = 63 AND Y = 9 else "111111110000" when X = 64 AND Y = 9 else "111111110000" when X = 65 AND Y = 9 else "111111110000" when X = 66 AND Y = 9 else "111111110000" when X = 67 AND Y = 9 else "111111110000" when X = 68 AND Y = 9 else "111111110000" when X = 0 AND Y = 10 else "111111110000" when X = 1 AND Y = 10 else "111111110000" when X = 2 AND Y = 10 else "111111110000" when X = 3 AND Y = 10 else "111111110000" when X = 4 AND Y = 10 else "111111110000" when X = 5 AND Y = 10 else "111111110000" when X = 6 AND Y = 10 else "111111110000" when X = 7 AND Y = 10 else "111111110000" when X = 8 AND Y = 10 else "010101110111" when X = 9 AND Y = 10 else "001100110011" when X = 10 AND Y = 10 else "100010001000" when X = 11 AND Y = 10 else "011101110111" when X = 12 AND Y = 10 else "000100010001" when X = 13 AND Y = 10 else "000000000000" when X = 14 AND Y = 10 else "000000000000" when X = 15 AND Y = 10 else "000100100010" when X = 16 AND Y = 10 else "100010111101" when X = 17 AND Y = 10 else "111111110000" when X = 18 AND Y = 10 else "100001101011" when X = 19 AND Y = 10 else "011100101001" when X = 20 AND Y = 10 else "011100101001" when X = 21 AND Y = 10 else "100100111000" when X = 22 AND Y = 10 else "111110000011" when X = 23 AND Y = 10 else "111110000000" when X = 24 AND Y = 10 else "111101000000" when X = 25 AND Y = 10 else "111100010000" when X = 26 AND Y = 10 else "101101100110" when X = 27 AND Y = 10 else "000010101101" when X = 28 AND Y = 10 else "000100011111" when X = 29 AND Y = 10 else "000100101111" when X = 30 AND Y = 10 else "101110110110" when X = 31 AND Y = 10 else "111111110000" when X = 32 AND Y = 10 else "111111110000" when X = 33 AND Y = 10 else "111111110000" when X = 34 AND Y = 10 else "110111010100" when X = 35 AND Y = 10 else "001000111110" when X = 36 AND Y = 10 else "000100001111" when X = 37 AND Y = 10 else "000010001110" when X = 38 AND Y = 10 else "100110001000" when X = 39 AND Y = 10 else "111100100001" when X = 40 AND Y = 10 else "111100010000" when X = 41 AND Y = 10 else "111101110000" when X = 42 AND Y = 10 else "111110010001" when X = 43 AND Y = 10 else "110001100110" when X = 44 AND Y = 10 else "011100101001" when X = 45 AND Y = 10 else "011100101001" when X = 46 AND Y = 10 else "011100101010" when X = 47 AND Y = 10 else "100110101101" when X = 48 AND Y = 10 else "111111110000" when X = 49 AND Y = 10 else "010101111000" when X = 50 AND Y = 10 else "000000000000" when X = 51 AND Y = 10 else "000000000000" when X = 52 AND Y = 10 else "000000000000" when X = 53 AND Y = 10 else "011001100110" when X = 54 AND Y = 10 else "100010001000" when X = 55 AND Y = 10 else "010001000100" when X = 56 AND Y = 10 else "001101010101" when X = 57 AND Y = 10 else "111111110000" when X = 58 AND Y = 10 else "111111110000" when X = 59 AND Y = 10 else "111111110000" when X = 60 AND Y = 10 else "111111110000" when X = 61 AND Y = 10 else "111111110000" when X = 62 AND Y = 10 else "111111110000" when X = 63 AND Y = 10 else "111111110000" when X = 64 AND Y = 10 else "111111110000" when X = 65 AND Y = 10 else "111111110000" when X = 66 AND Y = 10 else "111111110000" when X = 67 AND Y = 10 else "111111110000" when X = 68 AND Y = 10 else "111111110000" when X = 0 AND Y = 11 else "111111110000" when X = 1 AND Y = 11 else "111111110000" when X = 2 AND Y = 11 else "111111110000" when X = 3 AND Y = 11 else "111111110000" when X = 4 AND Y = 11 else "111111110000" when X = 5 AND Y = 11 else "111111110000" when X = 6 AND Y = 11 else "111111110000" when X = 7 AND Y = 11 else "111111110000" when X = 8 AND Y = 11 else "010001110111" when X = 9 AND Y = 11 else "000000000000" when X = 10 AND Y = 11 else "000100010001" when X = 11 AND Y = 11 else "000100010001" when X = 12 AND Y = 11 else "000000000000" when X = 13 AND Y = 11 else "000000000000" when X = 14 AND Y = 11 else "000000000000" when X = 15 AND Y = 11 else "000100000001" when X = 16 AND Y = 11 else "011100111001" when X = 17 AND Y = 11 else "011100111010" when X = 18 AND Y = 11 else "011100011010" when X = 19 AND Y = 11 else "101001000111" when X = 20 AND Y = 11 else "111001110011" when X = 21 AND Y = 11 else "111001110011" when X = 22 AND Y = 11 else "111110000000" when X = 23 AND Y = 11 else "111110000000" when X = 24 AND Y = 11 else "111100110000" when X = 25 AND Y = 11 else "101101110110" when X = 26 AND Y = 11 else "001110001100" when X = 27 AND Y = 11 else "000100101111" when X = 28 AND Y = 11 else "000100101111" when X = 29 AND Y = 11 else "101010110111" when X = 30 AND Y = 11 else "111011100010" when X = 31 AND Y = 11 else "111111110000" when X = 32 AND Y = 11 else "111111110000" when X = 33 AND Y = 11 else "111111110000" when X = 34 AND Y = 11 else "111011100001" when X = 35 AND Y = 11 else "110011000101" when X = 36 AND Y = 11 else "001001001101" when X = 37 AND Y = 11 else "000100011111" when X = 38 AND Y = 11 else "001001111101" when X = 39 AND Y = 11 else "011110101010" when X = 40 AND Y = 11 else "111000110010" when X = 41 AND Y = 11 else "111101110000" when X = 42 AND Y = 11 else "111110010000" when X = 43 AND Y = 11 else "111110000001" when X = 44 AND Y = 11 else "111001110011" when X = 45 AND Y = 11 else "110101100100" when X = 46 AND Y = 11 else "011100101001" when X = 47 AND Y = 11 else "011100111010" when X = 48 AND Y = 11 else "011100111010" when X = 49 AND Y = 11 else "010000100101" when X = 50 AND Y = 11 else "000000000000" when X = 51 AND Y = 11 else "000000000000" when X = 52 AND Y = 11 else "000000000000" when X = 53 AND Y = 11 else "000100010001" when X = 54 AND Y = 11 else "000100010001" when X = 55 AND Y = 11 else "000000000000" when X = 56 AND Y = 11 else "001101000100" when X = 57 AND Y = 11 else "111111110000" when X = 58 AND Y = 11 else "111111110000" when X = 59 AND Y = 11 else "111111110000" when X = 60 AND Y = 11 else "111111110000" when X = 61 AND Y = 11 else "111111110000" when X = 62 AND Y = 11 else "111111110000" when X = 63 AND Y = 11 else "111111110000" when X = 64 AND Y = 11 else "111111110000" when X = 65 AND Y = 11 else "111111110000" when X = 66 AND Y = 11 else "111111110000" when X = 67 AND Y = 11 else "111111110000" when X = 68 AND Y = 11 else "111111110000" when X = 0 AND Y = 12 else "111111110000" when X = 1 AND Y = 12 else "111111110000" when X = 2 AND Y = 12 else "111111110000" when X = 3 AND Y = 12 else "111111110000" when X = 4 AND Y = 12 else "111111110000" when X = 5 AND Y = 12 else "111111110000" when X = 6 AND Y = 12 else "111111110000" when X = 7 AND Y = 12 else "111111110000" when X = 8 AND Y = 12 else "010001110111" when X = 9 AND Y = 12 else "000000000000" when X = 10 AND Y = 12 else "000000000000" when X = 11 AND Y = 12 else "000000000000" when X = 12 AND Y = 12 else "000000000000" when X = 13 AND Y = 12 else "000000000000" when X = 14 AND Y = 12 else "001000010000" when X = 15 AND Y = 12 else "101001100001" when X = 16 AND Y = 12 else "110001100100" when X = 17 AND Y = 12 else "110101100100" when X = 18 AND Y = 12 else "110101100101" when X = 19 AND Y = 12 else "111001110011" when X = 20 AND Y = 12 else "111110010000" when X = 21 AND Y = 12 else "111110010000" when X = 22 AND Y = 12 else "111110000000" when X = 23 AND Y = 12 else "111110000000" when X = 24 AND Y = 12 else "111100110000" when X = 25 AND Y = 12 else "101010000111" when X = 26 AND Y = 12 else "000010011110" when X = 27 AND Y = 12 else "000100001111" when X = 28 AND Y = 12 else "000100101111" when X = 29 AND Y = 12 else "110111010100" when X = 30 AND Y = 12 else "111111110000" when X = 31 AND Y = 12 else "111111110000" when X = 32 AND Y = 12 else "111111110000" when X = 33 AND Y = 12 else "111111110000" when X = 34 AND Y = 12 else "111111110000" when X = 35 AND Y = 12 else "111011100010" when X = 36 AND Y = 12 else "001101001101" when X = 37 AND Y = 12 else "000100001111" when X = 38 AND Y = 12 else "000001101110" when X = 39 AND Y = 12 else "010011001100" when X = 40 AND Y = 12 else "111000110010" when X = 41 AND Y = 12 else "111101110000" when X = 42 AND Y = 12 else "111110010000" when X = 43 AND Y = 12 else "111110010000" when X = 44 AND Y = 12 else "111110010000" when X = 45 AND Y = 12 else "111110000001" when X = 46 AND Y = 12 else "110101100100" when X = 47 AND Y = 12 else "110101100100" when X = 48 AND Y = 12 else "110101100100" when X = 49 AND Y = 12 else "110001100011" when X = 50 AND Y = 12 else "011101000000" when X = 51 AND Y = 12 else "000000000000" when X = 52 AND Y = 12 else "000000000000" when X = 53 AND Y = 12 else "000000000000" when X = 54 AND Y = 12 else "000000000000" when X = 55 AND Y = 12 else "000000000000" when X = 56 AND Y = 12 else "001101000100" when X = 57 AND Y = 12 else "111111110000" when X = 58 AND Y = 12 else "111111110000" when X = 59 AND Y = 12 else "111111110000" when X = 60 AND Y = 12 else "111111110000" when X = 61 AND Y = 12 else "111111110000" when X = 62 AND Y = 12 else "111111110000" when X = 63 AND Y = 12 else "111111110000" when X = 64 AND Y = 12 else "111111110000" when X = 65 AND Y = 12 else "111111110000" when X = 66 AND Y = 12 else "111111110000" when X = 67 AND Y = 12 else "111111110000" when X = 68 AND Y = 12 else "111111110000" when X = 0 AND Y = 13 else "111111110000" when X = 1 AND Y = 13 else "111111110000" when X = 2 AND Y = 13 else "111111110000" when X = 3 AND Y = 13 else "111111110000" when X = 4 AND Y = 13 else "111111110000" when X = 5 AND Y = 13 else "111111110000" when X = 6 AND Y = 13 else "111111110000" when X = 7 AND Y = 13 else "111111110000" when X = 8 AND Y = 13 else "010001110111" when X = 9 AND Y = 13 else "000000000000" when X = 10 AND Y = 13 else "000000000000" when X = 11 AND Y = 13 else "000000000000" when X = 12 AND Y = 13 else "000000000000" when X = 13 AND Y = 13 else "001100010000" when X = 14 AND Y = 13 else "101001010000" when X = 15 AND Y = 13 else "111110010000" when X = 16 AND Y = 13 else "111110010000" when X = 17 AND Y = 13 else "111110010000" when X = 18 AND Y = 13 else "111110010000" when X = 19 AND Y = 13 else "111110010000" when X = 20 AND Y = 13 else "111110000000" when X = 21 AND Y = 13 else "111110000000" when X = 22 AND Y = 13 else "111110000000" when X = 23 AND Y = 13 else "111110010000" when X = 24 AND Y = 13 else "110010000101" when X = 25 AND Y = 13 else "011110101010" when X = 26 AND Y = 13 else "000010011110" when X = 27 AND Y = 13 else "001000011110" when X = 28 AND Y = 13 else "100001011001" when X = 29 AND Y = 13 else "111010110011" when X = 30 AND Y = 13 else "111111000000" when X = 31 AND Y = 13 else "111111000000" when X = 32 AND Y = 13 else "111111000000" when X = 33 AND Y = 13 else "111111000000" when X = 34 AND Y = 13 else "111111000000" when X = 35 AND Y = 13 else "111110110001" when X = 36 AND Y = 13 else "100101111000" when X = 37 AND Y = 13 else "001100101101" when X = 38 AND Y = 13 else "000001101111" when X = 39 AND Y = 13 else "001111001100" when X = 40 AND Y = 13 else "100110001000" when X = 41 AND Y = 13 else "111010000011" when X = 42 AND Y = 13 else "111110000000" when X = 43 AND Y = 13 else "111110000000" when X = 44 AND Y = 13 else "111110000000" when X = 45 AND Y = 13 else "111110000000" when X = 46 AND Y = 13 else "111110010000" when X = 47 AND Y = 13 else "111110010000" when X = 48 AND Y = 13 else "111110010000" when X = 49 AND Y = 13 else "111110010000" when X = 50 AND Y = 13 else "111001110000" when X = 51 AND Y = 13 else "011000110000" when X = 52 AND Y = 13 else "000000000000" when X = 53 AND Y = 13 else "000000000000" when X = 54 AND Y = 13 else "000000000000" when X = 55 AND Y = 13 else "000000000000" when X = 56 AND Y = 13 else "001101000100" when X = 57 AND Y = 13 else "111111110000" when X = 58 AND Y = 13 else "111111110000" when X = 59 AND Y = 13 else "111111110000" when X = 60 AND Y = 13 else "111111110000" when X = 61 AND Y = 13 else "111111110000" when X = 62 AND Y = 13 else "111111110000" when X = 63 AND Y = 13 else "111111110000" when X = 64 AND Y = 13 else "111111110000" when X = 65 AND Y = 13 else "111111110000" when X = 66 AND Y = 13 else "111111110000" when X = 67 AND Y = 13 else "111111110000" when X = 68 AND Y = 13 else "111111110000" when X = 0 AND Y = 14 else "111111110000" when X = 1 AND Y = 14 else "111111110000" when X = 2 AND Y = 14 else "111111110000" when X = 3 AND Y = 14 else "111111110000" when X = 4 AND Y = 14 else "111111110000" when X = 5 AND Y = 14 else "111111110000" when X = 6 AND Y = 14 else "111111110000" when X = 7 AND Y = 14 else "111111110000" when X = 8 AND Y = 14 else "010001110111" when X = 9 AND Y = 14 else "000000000000" when X = 10 AND Y = 14 else "000000000000" when X = 11 AND Y = 14 else "000000000000" when X = 12 AND Y = 14 else "010000100000" when X = 13 AND Y = 14 else "101001010000" when X = 14 AND Y = 14 else "111110010000" when X = 15 AND Y = 14 else "111110000000" when X = 16 AND Y = 14 else "111101110000" when X = 17 AND Y = 14 else "111110000000" when X = 18 AND Y = 14 else "111110010000" when X = 19 AND Y = 14 else "111110010000" when X = 20 AND Y = 14 else "111110010000" when X = 21 AND Y = 14 else "111110010000" when X = 22 AND Y = 14 else "111110010000" when X = 23 AND Y = 14 else "111110010000" when X = 24 AND Y = 14 else "011111001010" when X = 25 AND Y = 14 else "000011011101" when X = 26 AND Y = 14 else "001110011100" when X = 27 AND Y = 14 else "011101011010" when X = 28 AND Y = 14 else "111110000001" when X = 29 AND Y = 14 else "111110000000" when X = 30 AND Y = 14 else "111110000000" when X = 31 AND Y = 14 else "111110000000" when X = 32 AND Y = 14 else "111110000000" when X = 33 AND Y = 14 else "111110000000" when X = 34 AND Y = 14 else "111110000000" when X = 35 AND Y = 14 else "111110000000" when X = 36 AND Y = 14 else "111110010000" when X = 37 AND Y = 14 else "100101101000" when X = 38 AND Y = 14 else "010010001100" when X = 39 AND Y = 14 else "000011011101" when X = 40 AND Y = 14 else "000011011101" when X = 41 AND Y = 14 else "110010100101" when X = 42 AND Y = 14 else "111110000000" when X = 43 AND Y = 14 else "111110010000" when X = 44 AND Y = 14 else "111110010000" when X = 45 AND Y = 14 else "111110010000" when X = 46 AND Y = 14 else "111110010000" when X = 47 AND Y = 14 else "111110010000" when X = 48 AND Y = 14 else "111101110000" when X = 49 AND Y = 14 else "111101110000" when X = 50 AND Y = 14 else "111110010000" when X = 51 AND Y = 14 else "111010000000" when X = 52 AND Y = 14 else "010100110000" when X = 53 AND Y = 14 else "000000000000" when X = 54 AND Y = 14 else "000000000000" when X = 55 AND Y = 14 else "000000000000" when X = 56 AND Y = 14 else "001101000100" when X = 57 AND Y = 14 else "111111110000" when X = 58 AND Y = 14 else "111111110000" when X = 59 AND Y = 14 else "111111110000" when X = 60 AND Y = 14 else "111111110000" when X = 61 AND Y = 14 else "111111110000" when X = 62 AND Y = 14 else "111111110000" when X = 63 AND Y = 14 else "111111110000" when X = 64 AND Y = 14 else "111111110000" when X = 65 AND Y = 14 else "111111110000" when X = 66 AND Y = 14 else "111111110000" when X = 67 AND Y = 14 else "111111110000" when X = 68 AND Y = 14 else "111111110000" when X = 0 AND Y = 15 else "111111110000" when X = 1 AND Y = 15 else "111111110000" when X = 2 AND Y = 15 else "111111110000" when X = 3 AND Y = 15 else "111111110000" when X = 4 AND Y = 15 else "111111110000" when X = 5 AND Y = 15 else "111111110000" when X = 6 AND Y = 15 else "111111110000" when X = 7 AND Y = 15 else "111111110000" when X = 8 AND Y = 15 else "010001110111" when X = 9 AND Y = 15 else "000000000000" when X = 10 AND Y = 15 else "000000000000" when X = 11 AND Y = 15 else "001100100000" when X = 12 AND Y = 15 else "110101110000" when X = 13 AND Y = 15 else "111110010000" when X = 14 AND Y = 15 else "111110010000" when X = 15 AND Y = 15 else "111110000000" when X = 16 AND Y = 15 else "111100100000" when X = 17 AND Y = 15 else "111101100000" when X = 18 AND Y = 15 else "111101110000" when X = 19 AND Y = 15 else "111101110000" when X = 20 AND Y = 15 else "111101110000" when X = 21 AND Y = 15 else "111101110000" when X = 22 AND Y = 15 else "111101110000" when X = 23 AND Y = 15 else "111101110000" when X = 24 AND Y = 15 else "100110101000" when X = 25 AND Y = 15 else "010110111011" when X = 26 AND Y = 15 else "101010101000" when X = 27 AND Y = 15 else "111101110000" when X = 28 AND Y = 15 else "111101110000" when X = 29 AND Y = 15 else "111101110000" when X = 30 AND Y = 15 else "111101110000" when X = 31 AND Y = 15 else "111101110000" when X = 32 AND Y = 15 else "111101110000" when X = 33 AND Y = 15 else "111101110000" when X = 34 AND Y = 15 else "111101110000" when X = 35 AND Y = 15 else "111101110000" when X = 36 AND Y = 15 else "111101110000" when X = 37 AND Y = 15 else "111101110000" when X = 38 AND Y = 15 else "101110010110" when X = 39 AND Y = 15 else "011010111011" when X = 40 AND Y = 15 else "011010111011" when X = 41 AND Y = 15 else "110110000100" when X = 42 AND Y = 15 else "111101110000" when X = 43 AND Y = 15 else "111101110000" when X = 44 AND Y = 15 else "111101110000" when X = 45 AND Y = 15 else "111101110000" when X = 46 AND Y = 15 else "111101110000" when X = 47 AND Y = 15 else "111101110000" when X = 48 AND Y = 15 else "111100110000" when X = 49 AND Y = 15 else "111101010000" when X = 50 AND Y = 15 else "111110010000" when X = 51 AND Y = 15 else "111110000000" when X = 52 AND Y = 15 else "111110000000" when X = 53 AND Y = 15 else "010100110000" when X = 54 AND Y = 15 else "000000000000" when X = 55 AND Y = 15 else "000000000000" when X = 56 AND Y = 15 else "001101000100" when X = 57 AND Y = 15 else "111111110000" when X = 58 AND Y = 15 else "111111110000" when X = 59 AND Y = 15 else "111111110000" when X = 60 AND Y = 15 else "111111110000" when X = 61 AND Y = 15 else "111111110000" when X = 62 AND Y = 15 else "111111110000" when X = 63 AND Y = 15 else "111111110000" when X = 64 AND Y = 15 else "111111110000" when X = 65 AND Y = 15 else "111111110000" when X = 66 AND Y = 15 else "111111110000" when X = 67 AND Y = 15 else "111111110000" when X = 68 AND Y = 15 else "111111110000" when X = 0 AND Y = 16 else "111111110000" when X = 1 AND Y = 16 else "111111110000" when X = 2 AND Y = 16 else "111111110000" when X = 3 AND Y = 16 else "111111110000" when X = 4 AND Y = 16 else "111111110000" when X = 5 AND Y = 16 else "111111110000" when X = 6 AND Y = 16 else "111111110000" when X = 7 AND Y = 16 else "111111110000" when X = 8 AND Y = 16 else "010101110111" when X = 9 AND Y = 16 else "000000000000" when X = 10 AND Y = 16 else "001100100000" when X = 11 AND Y = 16 else "111001110000" when X = 12 AND Y = 16 else "111110000000" when X = 13 AND Y = 16 else "111110000000" when X = 14 AND Y = 16 else "111110010000" when X = 15 AND Y = 16 else "111110000000" when X = 16 AND Y = 16 else "111100010000" when X = 17 AND Y = 16 else "111100010000" when X = 18 AND Y = 16 else "111100010000" when X = 19 AND Y = 16 else "111100010000" when X = 20 AND Y = 16 else "111100010000" when X = 21 AND Y = 16 else "111100010000" when X = 22 AND Y = 16 else "111100010000" when X = 23 AND Y = 16 else "111100010000" when X = 24 AND Y = 16 else "111100100001" when X = 25 AND Y = 16 else "111000100001" when X = 26 AND Y = 16 else "111100100001" when X = 27 AND Y = 16 else "111100010000" when X = 28 AND Y = 16 else "111100010000" when X = 29 AND Y = 16 else "111100010000" when X = 30 AND Y = 16 else "111100010000" when X = 31 AND Y = 16 else "111100010000" when X = 32 AND Y = 16 else "111100010000" when X = 33 AND Y = 16 else "111100010000" when X = 34 AND Y = 16 else "111100010000" when X = 35 AND Y = 16 else "111100010000" when X = 36 AND Y = 16 else "111100010000" when X = 37 AND Y = 16 else "111100010000" when X = 38 AND Y = 16 else "111100010001" when X = 39 AND Y = 16 else "111000100001" when X = 40 AND Y = 16 else "111000100001" when X = 41 AND Y = 16 else "111100010000" when X = 42 AND Y = 16 else "111100010000" when X = 43 AND Y = 16 else "111100010000" when X = 44 AND Y = 16 else "111100010000" when X = 45 AND Y = 16 else "111100010000" when X = 46 AND Y = 16 else "111100010000" when X = 47 AND Y = 16 else "111100010000" when X = 48 AND Y = 16 else "111100000000" when X = 49 AND Y = 16 else "111101010000" when X = 50 AND Y = 16 else "111110010000" when X = 51 AND Y = 16 else "111110000000" when X = 52 AND Y = 16 else "111110000000" when X = 53 AND Y = 16 else "111110000000" when X = 54 AND Y = 16 else "010100110000" when X = 55 AND Y = 16 else "000000000000" when X = 56 AND Y = 16 else "010001000100" when X = 57 AND Y = 16 else "111111110000" when X = 58 AND Y = 16 else "111111110000" when X = 59 AND Y = 16 else "111111110000" when X = 60 AND Y = 16 else "111111110000" when X = 61 AND Y = 16 else "111111110000" when X = 62 AND Y = 16 else "111111110000" when X = 63 AND Y = 16 else "111111110000" when X = 64 AND Y = 16 else "111111110000" when X = 65 AND Y = 16 else "111111110000" when X = 66 AND Y = 16 else "111111110000" when X = 67 AND Y = 16 else "111111110000" when X = 68 AND Y = 16 else "111111110000" when X = 0 AND Y = 17 else "111111110000" when X = 1 AND Y = 17 else "111111110000" when X = 2 AND Y = 17 else "111111110000" when X = 3 AND Y = 17 else "111111110000" when X = 4 AND Y = 17 else "111111110000" when X = 5 AND Y = 17 else "111111110000" when X = 6 AND Y = 17 else "111111110000" when X = 7 AND Y = 17 else "110110111000" when X = 8 AND Y = 17 else "111010000010" when X = 9 AND Y = 17 else "110101110000" when X = 10 AND Y = 17 else "110101110000" when X = 11 AND Y = 17 else "111110000000" when X = 12 AND Y = 17 else "111110000000" when X = 13 AND Y = 17 else "111110000000" when X = 14 AND Y = 17 else "111110010000" when X = 15 AND Y = 17 else "111110000000" when X = 16 AND Y = 17 else "111100010000" when X = 17 AND Y = 17 else "101100000000" when X = 18 AND Y = 17 else "101000000000" when X = 19 AND Y = 17 else "101000000000" when X = 20 AND Y = 17 else "101000000000" when X = 21 AND Y = 17 else "101000000000" when X = 22 AND Y = 17 else "101000000000" when X = 23 AND Y = 17 else "101000000000" when X = 24 AND Y = 17 else "101000000000" when X = 25 AND Y = 17 else "101000000000" when X = 26 AND Y = 17 else "101000000000" when X = 27 AND Y = 17 else "101000000000" when X = 28 AND Y = 17 else "101000000000" when X = 29 AND Y = 17 else "101000000000" when X = 30 AND Y = 17 else "101000000000" when X = 31 AND Y = 17 else "101000000000" when X = 32 AND Y = 17 else "101000000000" when X = 33 AND Y = 17 else "101000000000" when X = 34 AND Y = 17 else "101000000000" when X = 35 AND Y = 17 else "101000000000" when X = 36 AND Y = 17 else "101000000000" when X = 37 AND Y = 17 else "101000000000" when X = 38 AND Y = 17 else "101000000000" when X = 39 AND Y = 17 else "101000000000" when X = 40 AND Y = 17 else "101000000000" when X = 41 AND Y = 17 else "101000000000" when X = 42 AND Y = 17 else "101000000000" when X = 43 AND Y = 17 else "101000000000" when X = 44 AND Y = 17 else "101000000000" when X = 45 AND Y = 17 else "101000000000" when X = 46 AND Y = 17 else "101000000000" when X = 47 AND Y = 17 else "101000000000" when X = 48 AND Y = 17 else "110100000000" when X = 49 AND Y = 17 else "111101010000" when X = 50 AND Y = 17 else "111110010000" when X = 51 AND Y = 17 else "111110000000" when X = 52 AND Y = 17 else "111110000000" when X = 53 AND Y = 17 else "111110000000" when X = 54 AND Y = 17 else "111001110000" when X = 55 AND Y = 17 else "110101110000" when X = 56 AND Y = 17 else "110110000001" when X = 57 AND Y = 17 else "110110100110" when X = 58 AND Y = 17 else "111111110000" when X = 59 AND Y = 17 else "111111110000" when X = 60 AND Y = 17 else "111111110000" when X = 61 AND Y = 17 else "111111110000" when X = 62 AND Y = 17 else "111111110000" when X = 63 AND Y = 17 else "111111110000" when X = 64 AND Y = 17 else "111111110000" when X = 65 AND Y = 17 else "111111110000" when X = 66 AND Y = 17 else "111111110000" when X = 67 AND Y = 17 else "111111110000" when X = 68 AND Y = 17 else "111111110000" when X = 0 AND Y = 18 else "111111110000" when X = 1 AND Y = 18 else "111111110000" when X = 2 AND Y = 18 else "011010011010" when X = 3 AND Y = 18 else "001101000100" when X = 4 AND Y = 18 else "001101000100" when X = 5 AND Y = 18 else "001101000100" when X = 6 AND Y = 18 else "001101000100" when X = 7 AND Y = 18 else "010000110010" when X = 8 AND Y = 18 else "010100100000" when X = 9 AND Y = 18 else "010100110000" when X = 10 AND Y = 18 else "010100110000" when X = 11 AND Y = 18 else "010100100000" when X = 12 AND Y = 18 else "010100100000" when X = 13 AND Y = 18 else "101001010000" when X = 14 AND Y = 18 else "111110010000" when X = 15 AND Y = 18 else "111110000000" when X = 16 AND Y = 18 else "111100010000" when X = 17 AND Y = 18 else "101000000000" when X = 18 AND Y = 18 else "100000000000" when X = 19 AND Y = 18 else "100000000000" when X = 20 AND Y = 18 else "100000000000" when X = 21 AND Y = 18 else "100000000000" when X = 22 AND Y = 18 else "100000000000" when X = 23 AND Y = 18 else "100000000000" when X = 24 AND Y = 18 else "100000000000" when X = 25 AND Y = 18 else "100000000000" when X = 26 AND Y = 18 else "100000000000" when X = 27 AND Y = 18 else "100000000000" when X = 28 AND Y = 18 else "100000000000" when X = 29 AND Y = 18 else "100000000000" when X = 30 AND Y = 18 else "100000000000" when X = 31 AND Y = 18 else "100000000000" when X = 32 AND Y = 18 else "100000000000" when X = 33 AND Y = 18 else "100000000000" when X = 34 AND Y = 18 else "100000000000" when X = 35 AND Y = 18 else "100000000000" when X = 36 AND Y = 18 else "100000000000" when X = 37 AND Y = 18 else "100000000000" when X = 38 AND Y = 18 else "100000000000" when X = 39 AND Y = 18 else "100000000000" when X = 40 AND Y = 18 else "100000000000" when X = 41 AND Y = 18 else "100000000000" when X = 42 AND Y = 18 else "100000000000" when X = 43 AND Y = 18 else "100000000000" when X = 44 AND Y = 18 else "100000000000" when X = 45 AND Y = 18 else "100000000000" when X = 46 AND Y = 18 else "100000000000" when X = 47 AND Y = 18 else "100000000000" when X = 48 AND Y = 18 else "110100000000" when X = 49 AND Y = 18 else "111101010000" when X = 50 AND Y = 18 else "111110010000" when X = 51 AND Y = 18 else "111010000000" when X = 52 AND Y = 18 else "011000110000" when X = 53 AND Y = 18 else "010100100000" when X = 54 AND Y = 18 else "010100110000" when X = 55 AND Y = 18 else "010100110000" when X = 56 AND Y = 18 else "010100110000" when X = 57 AND Y = 18 else "010000110001" when X = 58 AND Y = 18 else "001101000100" when X = 59 AND Y = 18 else "001101000100" when X = 60 AND Y = 18 else "001101000100" when X = 61 AND Y = 18 else "001101000100" when X = 62 AND Y = 18 else "010101111000" when X = 63 AND Y = 18 else "111111110000" when X = 64 AND Y = 18 else "111111110000" when X = 65 AND Y = 18 else "111111110000" when X = 66 AND Y = 18 else "111111110000" when X = 67 AND Y = 18 else "111111110000" when X = 68 AND Y = 18 else "111111110000" when X = 0 AND Y = 19 else "111111110000" when X = 1 AND Y = 19 else "100010111100" when X = 2 AND Y = 19 else "010001010110" when X = 3 AND Y = 19 else "000000000000" when X = 4 AND Y = 19 else "000000000000" when X = 5 AND Y = 19 else "000000000000" when X = 6 AND Y = 19 else "000000000000" when X = 7 AND Y = 19 else "000000000000" when X = 8 AND Y = 19 else "000000000000" when X = 9 AND Y = 19 else "000000000000" when X = 10 AND Y = 19 else "000000000000" when X = 11 AND Y = 19 else "000000000000" when X = 12 AND Y = 19 else "000000000000" when X = 13 AND Y = 19 else "010100100000" when X = 14 AND Y = 19 else "110101110000" when X = 15 AND Y = 19 else "111110000000" when X = 16 AND Y = 19 else "111100010000" when X = 17 AND Y = 19 else "101000000000" when X = 18 AND Y = 19 else "100000000000" when X = 19 AND Y = 19 else "100000000000" when X = 20 AND Y = 19 else "100000000000" when X = 21 AND Y = 19 else "100000000000" when X = 22 AND Y = 19 else "100000000000" when X = 23 AND Y = 19 else "100000000000" when X = 24 AND Y = 19 else "100000000000" when X = 25 AND Y = 19 else "100000000000" when X = 26 AND Y = 19 else "100000000000" when X = 27 AND Y = 19 else "100000000000" when X = 28 AND Y = 19 else "100000000000" when X = 29 AND Y = 19 else "100000000000" when X = 30 AND Y = 19 else "100000000000" when X = 31 AND Y = 19 else "100100000000" when X = 32 AND Y = 19 else "101000000000" when X = 33 AND Y = 19 else "101000000000" when X = 34 AND Y = 19 else "100100000000" when X = 35 AND Y = 19 else "100000000000" when X = 36 AND Y = 19 else "100000000000" when X = 37 AND Y = 19 else "100000000000" when X = 38 AND Y = 19 else "100000000000" when X = 39 AND Y = 19 else "100000000000" when X = 40 AND Y = 19 else "100000000000" when X = 41 AND Y = 19 else "100000000000" when X = 42 AND Y = 19 else "100000000000" when X = 43 AND Y = 19 else "100000000000" when X = 44 AND Y = 19 else "100000000000" when X = 45 AND Y = 19 else "100000000000" when X = 46 AND Y = 19 else "100000000000" when X = 47 AND Y = 19 else "100000000000" when X = 48 AND Y = 19 else "110100000000" when X = 49 AND Y = 19 else "111101010000" when X = 50 AND Y = 19 else "111110000000" when X = 51 AND Y = 19 else "101001010000" when X = 52 AND Y = 19 else "000100000000" when X = 53 AND Y = 19 else "000000000000" when X = 54 AND Y = 19 else "000000000000" when X = 55 AND Y = 19 else "000000000000" when X = 56 AND Y = 19 else "000000000000" when X = 57 AND Y = 19 else "000000000000" when X = 58 AND Y = 19 else "000000000000" when X = 59 AND Y = 19 else "000000000000" when X = 60 AND Y = 19 else "000000000000" when X = 61 AND Y = 19 else "000000000000" when X = 62 AND Y = 19 else "001000110100" when X = 63 AND Y = 19 else "011110111011" when X = 64 AND Y = 19 else "111111110000" when X = 65 AND Y = 19 else "111111110000" when X = 66 AND Y = 19 else "111111110000" when X = 67 AND Y = 19 else "111111110000" when X = 68 AND Y = 19 else "111111110000" when X = 0 AND Y = 20 else "111111110000" when X = 1 AND Y = 20 else "001101010110" when X = 2 AND Y = 20 else "000000000000" when X = 3 AND Y = 20 else "000000000000" when X = 4 AND Y = 20 else "000100010001" when X = 5 AND Y = 20 else "000100010001" when X = 6 AND Y = 20 else "000000000000" when X = 7 AND Y = 20 else "000000000000" when X = 8 AND Y = 20 else "000100010001" when X = 9 AND Y = 20 else "000100010001" when X = 10 AND Y = 20 else "000100010001" when X = 11 AND Y = 20 else "000100010001" when X = 12 AND Y = 20 else "000000000000" when X = 13 AND Y = 20 else "000000000000" when X = 14 AND Y = 20 else "010000100001" when X = 15 AND Y = 20 else "111001110011" when X = 16 AND Y = 20 else "111100010000" when X = 17 AND Y = 20 else "101000000000" when X = 18 AND Y = 20 else "100000000000" when X = 19 AND Y = 20 else "100000000000" when X = 20 AND Y = 20 else "100000000000" when X = 21 AND Y = 20 else "100000000000" when X = 22 AND Y = 20 else "100000000000" when X = 23 AND Y = 20 else "100000000000" when X = 24 AND Y = 20 else "100000000000" when X = 25 AND Y = 20 else "100000000000" when X = 26 AND Y = 20 else "100000000000" when X = 27 AND Y = 20 else "100000000000" when X = 28 AND Y = 20 else "100000000000" when X = 29 AND Y = 20 else "100000000000" when X = 30 AND Y = 20 else "100000000000" when X = 31 AND Y = 20 else "110000000000" when X = 32 AND Y = 20 else "111100000000" when X = 33 AND Y = 20 else "111000000000" when X = 34 AND Y = 20 else "100100000000" when X = 35 AND Y = 20 else "100000000000" when X = 36 AND Y = 20 else "100000000000" when X = 37 AND Y = 20 else "100000000000" when X = 38 AND Y = 20 else "100000000000" when X = 39 AND Y = 20 else "100000000000" when X = 40 AND Y = 20 else "100000000000" when X = 41 AND Y = 20 else "100000000000" when X = 42 AND Y = 20 else "100000000000" when X = 43 AND Y = 20 else "100000000000" when X = 44 AND Y = 20 else "100000000000" when X = 45 AND Y = 20 else "100000000000" when X = 46 AND Y = 20 else "100000000000" when X = 47 AND Y = 20 else "100000000000" when X = 48 AND Y = 20 else "110100000000" when X = 49 AND Y = 20 else "111101000010" when X = 50 AND Y = 20 else "101001100010" when X = 51 AND Y = 20 else "000000000000" when X = 52 AND Y = 20 else "000000000000" when X = 53 AND Y = 20 else "000000000000" when X = 54 AND Y = 20 else "000100010001" when X = 55 AND Y = 20 else "000100010001" when X = 56 AND Y = 20 else "000100010001" when X = 57 AND Y = 20 else "000000000000" when X = 58 AND Y = 20 else "000000000000" when X = 59 AND Y = 20 else "000000000000" when X = 60 AND Y = 20 else "000100010001" when X = 61 AND Y = 20 else "000000000000" when X = 62 AND Y = 20 else "000000000000" when X = 63 AND Y = 20 else "001000110011" when X = 64 AND Y = 20 else "111111110000" when X = 65 AND Y = 20 else "111111110000" when X = 66 AND Y = 20 else "111111110000" when X = 67 AND Y = 20 else "111111110000" when X = 68 AND Y = 20 else "111111110000" when X = 0 AND Y = 21 else "111111110000" when X = 1 AND Y = 21 else "001101010101" when X = 2 AND Y = 21 else "000000000000" when X = 3 AND Y = 21 else "001000100010" when X = 4 AND Y = 21 else "100010001000" when X = 5 AND Y = 21 else "011101110111" when X = 6 AND Y = 21 else "000100010001" when X = 7 AND Y = 21 else "010101010101" when X = 8 AND Y = 21 else "100010001000" when X = 9 AND Y = 21 else "100010001000" when X = 10 AND Y = 21 else "100010001000" when X = 11 AND Y = 21 else "011101110111" when X = 12 AND Y = 21 else "000100010001" when X = 13 AND Y = 21 else "000000000000" when X = 14 AND Y = 21 else "000000000100" when X = 15 AND Y = 21 else "001100101100" when X = 16 AND Y = 21 else "111000010010" when X = 17 AND Y = 21 else "101000000000" when X = 18 AND Y = 21 else "100000000000" when X = 19 AND Y = 21 else "100000000000" when X = 20 AND Y = 21 else "100000000000" when X = 21 AND Y = 21 else "100000000000" when X = 22 AND Y = 21 else "100000000000" when X = 23 AND Y = 21 else "100000000000" when X = 24 AND Y = 21 else "100000000000" when X = 25 AND Y = 21 else "100000000000" when X = 26 AND Y = 21 else "100000000000" when X = 27 AND Y = 21 else "100000000000" when X = 28 AND Y = 21 else "100000000000" when X = 29 AND Y = 21 else "100000000000" when X = 30 AND Y = 21 else "100000000000" when X = 31 AND Y = 21 else "110100000000" when X = 32 AND Y = 21 else "111100000000" when X = 33 AND Y = 21 else "111000000000" when X = 34 AND Y = 21 else "100100000000" when X = 35 AND Y = 21 else "100000000000" when X = 36 AND Y = 21 else "100000000000" when X = 37 AND Y = 21 else "100000000000" when X = 38 AND Y = 21 else "100000000000" when X = 39 AND Y = 21 else "100000000000" when X = 40 AND Y = 21 else "100000000000" when X = 41 AND Y = 21 else "100000000000" when X = 42 AND Y = 21 else "100000000000" when X = 43 AND Y = 21 else "100000000000" when X = 44 AND Y = 21 else "100000000000" when X = 45 AND Y = 21 else "100000000000" when X = 46 AND Y = 21 else "100000000000" when X = 47 AND Y = 21 else "100000000000" when X = 48 AND Y = 21 else "110100000000" when X = 49 AND Y = 21 else "100100100111" when X = 50 AND Y = 21 else "000100011010" when X = 51 AND Y = 21 else "000000000000" when X = 52 AND Y = 21 else "000000000000" when X = 53 AND Y = 21 else "011001100110" when X = 54 AND Y = 21 else "100010001000" when X = 55 AND Y = 21 else "100010001000" when X = 56 AND Y = 21 else "100010001000" when X = 57 AND Y = 21 else "011001100110" when X = 58 AND Y = 21 else "000100010001" when X = 59 AND Y = 21 else "011101110111" when X = 60 AND Y = 21 else "100010001000" when X = 61 AND Y = 21 else "001100110011" when X = 62 AND Y = 21 else "000000000000" when X = 63 AND Y = 21 else "001000100011" when X = 64 AND Y = 21 else "111111110000" when X = 65 AND Y = 21 else "111111110000" when X = 66 AND Y = 21 else "111111110000" when X = 67 AND Y = 21 else "111111110000" when X = 68 AND Y = 21 else "111111110000" when X = 0 AND Y = 22 else "111111110000" when X = 1 AND Y = 22 else "001101010101" when X = 2 AND Y = 22 else "000000000000" when X = 3 AND Y = 22 else "000000000000" when X = 4 AND Y = 22 else "001000100010" when X = 5 AND Y = 22 else "001000100010" when X = 6 AND Y = 22 else "000000000000" when X = 7 AND Y = 22 else "000100010001" when X = 8 AND Y = 22 else "001000100010" when X = 9 AND Y = 22 else "001000100010" when X = 10 AND Y = 22 else "001000100010" when X = 11 AND Y = 22 else "001000100010" when X = 12 AND Y = 22 else "000000000000" when X = 13 AND Y = 22 else "000000000000" when X = 14 AND Y = 22 else "000000000100" when X = 15 AND Y = 22 else "001000001101" when X = 16 AND Y = 22 else "110100010011" when X = 17 AND Y = 22 else "010100011010" when X = 18 AND Y = 22 else "001000001100" when X = 19 AND Y = 22 else "001000001100" when X = 20 AND Y = 22 else "001000001100" when X = 21 AND Y = 22 else "001000001100" when X = 22 AND Y = 22 else "001000001100" when X = 23 AND Y = 22 else "001000001100" when X = 24 AND Y = 22 else "001000001100" when X = 25 AND Y = 22 else "001000001100" when X = 26 AND Y = 22 else "001000001100" when X = 27 AND Y = 22 else "001000001100" when X = 28 AND Y = 22 else "001000001100" when X = 29 AND Y = 22 else "001000011100" when X = 30 AND Y = 22 else "101100010100" when X = 31 AND Y = 22 else "111100000000" when X = 32 AND Y = 22 else "111100000000" when X = 33 AND Y = 22 else "111100000000" when X = 34 AND Y = 22 else "110000000010" when X = 35 AND Y = 22 else "001100011011" when X = 36 AND Y = 22 else "001000001100" when X = 37 AND Y = 22 else "001000001100" when X = 38 AND Y = 22 else "001000001100" when X = 39 AND Y = 22 else "001000001100" when X = 40 AND Y = 22 else "001000001100" when X = 41 AND Y = 22 else "001000001100" when X = 42 AND Y = 22 else "001000001100" when X = 43 AND Y = 22 else "001000001100" when X = 44 AND Y = 22 else "001000001100" when X = 45 AND Y = 22 else "001000001100" when X = 46 AND Y = 22 else "001000001100" when X = 47 AND Y = 22 else "001000001100" when X = 48 AND Y = 22 else "101000010101" when X = 49 AND Y = 22 else "100100011000" when X = 50 AND Y = 22 else "000000001011" when X = 51 AND Y = 22 else "000000000000" when X = 52 AND Y = 22 else "000000000000" when X = 53 AND Y = 22 else "001000100010" when X = 54 AND Y = 22 else "001000100010" when X = 55 AND Y = 22 else "001000100010" when X = 56 AND Y = 22 else "001000100010" when X = 57 AND Y = 22 else "001000100010" when X = 58 AND Y = 22 else "000000000000" when X = 59 AND Y = 22 else "001000100010" when X = 60 AND Y = 22 else "001000100010" when X = 61 AND Y = 22 else "000100010001" when X = 62 AND Y = 22 else "000000000000" when X = 63 AND Y = 22 else "001000100011" when X = 64 AND Y = 22 else "111111110000" when X = 65 AND Y = 22 else "111111110000" when X = 66 AND Y = 22 else "111111110000" when X = 67 AND Y = 22 else "111111110000" when X = 68 AND Y = 22 else "111111110000" when X = 0 AND Y = 23 else "111111110000" when X = 1 AND Y = 23 else "001101010101" when X = 2 AND Y = 23 else "000000000000" when X = 3 AND Y = 23 else "000000000000" when X = 4 AND Y = 23 else "000000000000" when X = 5 AND Y = 23 else "000000000000" when X = 6 AND Y = 23 else "000000000000" when X = 7 AND Y = 23 else "000000000000" when X = 8 AND Y = 23 else "000000000000" when X = 9 AND Y = 23 else "000000000000" when X = 10 AND Y = 23 else "000000000000" when X = 11 AND Y = 23 else "000000000000" when X = 12 AND Y = 23 else "000000000000" when X = 13 AND Y = 23 else "000000000000" when X = 14 AND Y = 23 else "000000000100" when X = 15 AND Y = 23 else "001000011101" when X = 16 AND Y = 23 else "110100010011" when X = 17 AND Y = 23 else "001100011101" when X = 18 AND Y = 23 else "000100001111" when X = 19 AND Y = 23 else "000000111110" when X = 20 AND Y = 23 else "000001101100" when X = 21 AND Y = 23 else "000001101100" when X = 22 AND Y = 23 else "000001101100" when X = 23 AND Y = 23 else "000001101100" when X = 24 AND Y = 23 else "001100101100" when X = 25 AND Y = 23 else "010000001100" when X = 26 AND Y = 23 else "001100111100" when X = 27 AND Y = 23 else "000101011100" when X = 28 AND Y = 23 else "010000011100" when X = 29 AND Y = 23 else "010000001100" when X = 30 AND Y = 23 else "110000010100" when X = 31 AND Y = 23 else "111100000000" when X = 32 AND Y = 23 else "111100000000" when X = 33 AND Y = 23 else "111100000000" when X = 34 AND Y = 23 else "111000000010" when X = 35 AND Y = 23 else "010100011011" when X = 36 AND Y = 23 else "010000001100" when X = 37 AND Y = 23 else "001001001100" when X = 38 AND Y = 23 else "001001001100" when X = 39 AND Y = 23 else "010000001100" when X = 40 AND Y = 23 else "010000011100" when X = 41 AND Y = 23 else "000101001100" when X = 42 AND Y = 23 else "000001101100" when X = 43 AND Y = 23 else "000001101100" when X = 44 AND Y = 23 else "000001101100" when X = 45 AND Y = 23 else "000001011100" when X = 46 AND Y = 23 else "000100011111" when X = 47 AND Y = 23 else "000100001111" when X = 48 AND Y = 23 else "101000010111" when X = 49 AND Y = 23 else "100100011000" when X = 50 AND Y = 23 else "000000001011" when X = 51 AND Y = 23 else "000000000000" when X = 52 AND Y = 23 else "000000000000" when X = 53 AND Y = 23 else "000000000000" when X = 54 AND Y = 23 else "000000000000" when X = 55 AND Y = 23 else "000000000000" when X = 56 AND Y = 23 else "000000000000" when X = 57 AND Y = 23 else "000000000000" when X = 58 AND Y = 23 else "000000000000" when X = 59 AND Y = 23 else "000000000000" when X = 60 AND Y = 23 else "000000000000" when X = 61 AND Y = 23 else "000000000000" when X = 62 AND Y = 23 else "000000000000" when X = 63 AND Y = 23 else "001000100011" when X = 64 AND Y = 23 else "111111110000" when X = 65 AND Y = 23 else "111111110000" when X = 66 AND Y = 23 else "111111110000" when X = 67 AND Y = 23 else "111111110000" when X = 68 AND Y = 23 else "111111110000" when X = 0 AND Y = 24 else "111111110000" when X = 1 AND Y = 24 else "001101010101" when X = 2 AND Y = 24 else "000000000000" when X = 3 AND Y = 24 else "000000000000" when X = 4 AND Y = 24 else "000000000000" when X = 5 AND Y = 24 else "000000000000" when X = 6 AND Y = 24 else "000000000000" when X = 7 AND Y = 24 else "000000000000" when X = 8 AND Y = 24 else "000000000000" when X = 9 AND Y = 24 else "000000000000" when X = 10 AND Y = 24 else "000000000000" when X = 11 AND Y = 24 else "000000000000" when X = 12 AND Y = 24 else "000000000000" when X = 13 AND Y = 24 else "000000000000" when X = 14 AND Y = 24 else "000000000011" when X = 15 AND Y = 24 else "001100011100" when X = 16 AND Y = 24 else "100000011000" when X = 17 AND Y = 24 else "001000001110" when X = 18 AND Y = 24 else "000100001111" when X = 19 AND Y = 24 else "000001011100" when X = 20 AND Y = 24 else "000010011000" when X = 21 AND Y = 24 else "000010011000" when X = 22 AND Y = 24 else "000010001000" when X = 23 AND Y = 24 else "010001101001" when X = 24 AND Y = 24 else "011000101001" when X = 25 AND Y = 24 else "011100001001" when X = 26 AND Y = 24 else "010101001001" when X = 27 AND Y = 24 else "001101111001" when X = 28 AND Y = 24 else "011100011001" when X = 29 AND Y = 24 else "011100001001" when X = 30 AND Y = 24 else "110100000011" when X = 31 AND Y = 24 else "111100000000" when X = 32 AND Y = 24 else "111100000000" when X = 33 AND Y = 24 else "111100000000" when X = 34 AND Y = 24 else "111000000010" when X = 35 AND Y = 24 else "100000001000" when X = 36 AND Y = 24 else "011100001001" when X = 37 AND Y = 24 else "010001101001" when X = 38 AND Y = 24 else "010001011001" when X = 39 AND Y = 24 else "011100001001" when X = 40 AND Y = 24 else "011100011001" when X = 41 AND Y = 24 else "010101001001" when X = 42 AND Y = 24 else "001001111001" when X = 43 AND Y = 24 else "000010011000" when X = 44 AND Y = 24 else "000010011000" when X = 45 AND Y = 24 else "000010001001" when X = 46 AND Y = 24 else "000100011111" when X = 47 AND Y = 24 else "000100001111" when X = 48 AND Y = 24 else "010100011010" when X = 49 AND Y = 24 else "011000011010" when X = 50 AND Y = 24 else "001000001001" when X = 51 AND Y = 24 else "000000000000" when X = 52 AND Y = 24 else "000000000000" when X = 53 AND Y = 24 else "000000000000" when X = 54 AND Y = 24 else "000000000000" when X = 55 AND Y = 24 else "000000000000" when X = 56 AND Y = 24 else "000000000000" when X = 57 AND Y = 24 else "000000000000" when X = 58 AND Y = 24 else "000000000000" when X = 59 AND Y = 24 else "000000000000" when X = 60 AND Y = 24 else "000000000000" when X = 61 AND Y = 24 else "000000000000" when X = 62 AND Y = 24 else "000000000000" when X = 63 AND Y = 24 else "001000100011" when X = 64 AND Y = 24 else "111111110000" when X = 65 AND Y = 24 else "111111110000" when X = 66 AND Y = 24 else "111111110000" when X = 67 AND Y = 24 else "111111110000" when X = 68 AND Y = 24 else "111111110000" when X = 0 AND Y = 25 else "111111110000" when X = 1 AND Y = 25 else "001101010101" when X = 2 AND Y = 25 else "000000000000" when X = 3 AND Y = 25 else "000000000000" when X = 4 AND Y = 25 else "000000000000" when X = 5 AND Y = 25 else "000000000000" when X = 6 AND Y = 25 else "000000000000" when X = 7 AND Y = 25 else "000000000000" when X = 8 AND Y = 25 else "000000000000" when X = 9 AND Y = 25 else "000000000000" when X = 10 AND Y = 25 else "000000000000" when X = 11 AND Y = 25 else "000000000000" when X = 12 AND Y = 25 else "000000000000" when X = 13 AND Y = 25 else "000000000000" when X = 14 AND Y = 25 else "001000000010" when X = 15 AND Y = 25 else "011000001010" when X = 16 AND Y = 25 else "001000001110" when X = 17 AND Y = 25 else "000100001111" when X = 18 AND Y = 25 else "000100101111" when X = 19 AND Y = 25 else "000001101011" when X = 20 AND Y = 25 else "000010011000" when X = 21 AND Y = 25 else "000010011000" when X = 22 AND Y = 25 else "000110001001" when X = 23 AND Y = 25 else "011000101001" when X = 24 AND Y = 25 else "011100001001" when X = 25 AND Y = 25 else "011100001001" when X = 26 AND Y = 25 else "010101001001" when X = 27 AND Y = 25 else "001101111001" when X = 28 AND Y = 25 else "011000011001" when X = 29 AND Y = 25 else "011100001001" when X = 30 AND Y = 25 else "110100000011" when X = 31 AND Y = 25 else "111100000000" when X = 32 AND Y = 25 else "111100000000" when X = 33 AND Y = 25 else "111100000000" when X = 34 AND Y = 25 else "111000000010" when X = 35 AND Y = 25 else "011100001000" when X = 36 AND Y = 25 else "011000001001" when X = 37 AND Y = 25 else "010001101001" when X = 38 AND Y = 25 else "010001011001" when X = 39 AND Y = 25 else "011100001001" when X = 40 AND Y = 25 else "011100001001" when X = 41 AND Y = 25 else "011100001001" when X = 42 AND Y = 25 else "010001011001" when X = 43 AND Y = 25 else "000010011000" when X = 44 AND Y = 25 else "000010011000" when X = 45 AND Y = 25 else "000010001001" when X = 46 AND Y = 25 else "000000111101" when X = 47 AND Y = 25 else "000100011111" when X = 48 AND Y = 25 else "000100001111" when X = 49 AND Y = 25 else "010000001100" when X = 50 AND Y = 25 else "010100000110" when X = 51 AND Y = 25 else "000000000000" when X = 52 AND Y = 25 else "000000000000" when X = 53 AND Y = 25 else "000000000000" when X = 54 AND Y = 25 else "000000000000" when X = 55 AND Y = 25 else "000000000000" when X = 56 AND Y = 25 else "000000000000" when X = 57 AND Y = 25 else "000000000000" when X = 58 AND Y = 25 else "000000000000" when X = 59 AND Y = 25 else "000000000000" when X = 60 AND Y = 25 else "000000000000" when X = 61 AND Y = 25 else "000000000000" when X = 62 AND Y = 25 else "000000000000" when X = 63 AND Y = 25 else "001000100011" when X = 64 AND Y = 25 else "111111110000" when X = 65 AND Y = 25 else "111111110000" when X = 66 AND Y = 25 else "111111110000" when X = 67 AND Y = 25 else "111111110000" when X = 68 AND Y = 25 else "111111110000" when X = 0 AND Y = 26 else "111111110000" when X = 1 AND Y = 26 else "001101010101" when X = 2 AND Y = 26 else "000000000000" when X = 3 AND Y = 26 else "000000000000" when X = 4 AND Y = 26 else "000000000000" when X = 5 AND Y = 26 else "000000000000" when X = 6 AND Y = 26 else "000000000000" when X = 7 AND Y = 26 else "000000000000" when X = 8 AND Y = 26 else "000000000000" when X = 9 AND Y = 26 else "000000000000" when X = 10 AND Y = 26 else "000000000000" when X = 11 AND Y = 26 else "000000000000" when X = 12 AND Y = 26 else "000000000000" when X = 13 AND Y = 26 else "000000000000" when X = 14 AND Y = 26 else "000100000010" when X = 15 AND Y = 26 else "011000001001" when X = 16 AND Y = 26 else "011000001010" when X = 17 AND Y = 26 else "001000001110" when X = 18 AND Y = 26 else "000101011011" when X = 19 AND Y = 26 else "001010001001" when X = 20 AND Y = 26 else "001010001001" when X = 21 AND Y = 26 else "001010001001" when X = 22 AND Y = 26 else "001101111001" when X = 23 AND Y = 26 else "011000101001" when X = 24 AND Y = 26 else "011100001001" when X = 25 AND Y = 26 else "011100001001" when X = 26 AND Y = 26 else "010101001001" when X = 27 AND Y = 26 else "001101111001" when X = 28 AND Y = 26 else "011100101001" when X = 29 AND Y = 26 else "011100101001" when X = 30 AND Y = 26 else "110100100100" when X = 31 AND Y = 26 else "111100100001" when X = 32 AND Y = 26 else "111100100010" when X = 33 AND Y = 26 else "111100100001" when X = 34 AND Y = 26 else "111000100011" when X = 35 AND Y = 26 else "100000101001" when X = 36 AND Y = 26 else "011100101001" when X = 37 AND Y = 26 else "010001101001" when X = 38 AND Y = 26 else "010001011001" when X = 39 AND Y = 26 else "011100001001" when X = 40 AND Y = 26 else "011100001001" when X = 41 AND Y = 26 else "011100001001" when X = 42 AND Y = 26 else "010101011001" when X = 43 AND Y = 26 else "001010001001" when X = 44 AND Y = 26 else "001010001001" when X = 45 AND Y = 26 else "001010001001" when X = 46 AND Y = 26 else "001001111001" when X = 47 AND Y = 26 else "000100101101" when X = 48 AND Y = 26 else "010000001100" when X = 49 AND Y = 26 else "011100001010" when X = 50 AND Y = 26 else "010100000111" when X = 51 AND Y = 26 else "000000000000" when X = 52 AND Y = 26 else "000000000000" when X = 53 AND Y = 26 else "000000000000" when X = 54 AND Y = 26 else "000000000000" when X = 55 AND Y = 26 else "000000000000" when X = 56 AND Y = 26 else "000000000000" when X = 57 AND Y = 26 else "000000000000" when X = 58 AND Y = 26 else "000000000000" when X = 59 AND Y = 26 else "000000000000" when X = 60 AND Y = 26 else "000000000000" when X = 61 AND Y = 26 else "000000000000" when X = 62 AND Y = 26 else "000000000000" when X = 63 AND Y = 26 else "001000100011" when X = 64 AND Y = 26 else "111111110000" when X = 65 AND Y = 26 else "111111110000" when X = 66 AND Y = 26 else "111111110000" when X = 67 AND Y = 26 else "111111110000" when X = 68 AND Y = 26 else "111111110000" when X = 0 AND Y = 27 else "111111110000" when X = 1 AND Y = 27 else "001101010101" when X = 2 AND Y = 27 else "000000000000" when X = 3 AND Y = 27 else "000000000000" when X = 4 AND Y = 27 else "000000000000" when X = 5 AND Y = 27 else "000000000000" when X = 6 AND Y = 27 else "000000000000" when X = 7 AND Y = 27 else "000000000000" when X = 8 AND Y = 27 else "000000000000" when X = 9 AND Y = 27 else "000000000000" when X = 10 AND Y = 27 else "000000000000" when X = 11 AND Y = 27 else "000000000000" when X = 12 AND Y = 27 else "000000000000" when X = 13 AND Y = 27 else "000000000000" when X = 14 AND Y = 27 else "000100000010" when X = 15 AND Y = 27 else "011000001001" when X = 16 AND Y = 27 else "011100001001" when X = 17 AND Y = 27 else "011000001010" when X = 18 AND Y = 27 else "011000011010" when X = 19 AND Y = 27 else "011000101001" when X = 20 AND Y = 27 else "011000101001" when X = 21 AND Y = 27 else "011000101001" when X = 22 AND Y = 27 else "011000101001" when X = 23 AND Y = 27 else "011000011001" when X = 24 AND Y = 27 else "011100001001" when X = 25 AND Y = 27 else "011100001001" when X = 26 AND Y = 27 else "010101001001" when X = 27 AND Y = 27 else "001110001001" when X = 28 AND Y = 27 else "100110001001" when X = 29 AND Y = 27 else "100110001001" when X = 30 AND Y = 27 else "101010001001" when X = 31 AND Y = 27 else "101010011000" when X = 32 AND Y = 27 else "101010011000" when X = 33 AND Y = 27 else "101010011000" when X = 34 AND Y = 27 else "101010001001" when X = 35 AND Y = 27 else "100110001001" when X = 36 AND Y = 27 else "100110001001" when X = 37 AND Y = 27 else "010010011001" when X = 38 AND Y = 27 else "010001011001" when X = 39 AND Y = 27 else "011100001001" when X = 40 AND Y = 27 else "011100001001" when X = 41 AND Y = 27 else "011100001001" when X = 42 AND Y = 27 else "011000011001" when X = 43 AND Y = 27 else "011000101001" when X = 44 AND Y = 27 else "011000101001" when X = 45 AND Y = 27 else "011000101001" when X = 46 AND Y = 27 else "011000101001" when X = 47 AND Y = 27 else "011000011010" when X = 48 AND Y = 27 else "011000001010" when X = 49 AND Y = 27 else "011100001001" when X = 50 AND Y = 27 else "010100000111" when X = 51 AND Y = 27 else "000000000000" when X = 52 AND Y = 27 else "000000000000" when X = 53 AND Y = 27 else "000000000000" when X = 54 AND Y = 27 else "000000000000" when X = 55 AND Y = 27 else "000000000000" when X = 56 AND Y = 27 else "000000000000" when X = 57 AND Y = 27 else "000000000000" when X = 58 AND Y = 27 else "000000000000" when X = 59 AND Y = 27 else "000000000000" when X = 60 AND Y = 27 else "000000000000" when X = 61 AND Y = 27 else "000000000000" when X = 62 AND Y = 27 else "000000000000" when X = 63 AND Y = 27 else "001000110011" when X = 64 AND Y = 27 else "111111110000" when X = 65 AND Y = 27 else "111111110000" when X = 66 AND Y = 27 else "111111110000" when X = 67 AND Y = 27 else "111111110000" when X = 68 AND Y = 27 else "111111110000" when X = 0 AND Y = 28 else "111111110000" when X = 1 AND Y = 28 else "100010101010" when X = 2 AND Y = 28 else "010001000100" when X = 3 AND Y = 28 else "000000000000" when X = 4 AND Y = 28 else "000000000000" when X = 5 AND Y = 28 else "000000000000" when X = 6 AND Y = 28 else "000000000000" when X = 7 AND Y = 28 else "000000000000" when X = 8 AND Y = 28 else "000000000000" when X = 9 AND Y = 28 else "000000000000" when X = 10 AND Y = 28 else "000000000000" when X = 11 AND Y = 28 else "000000000000" when X = 12 AND Y = 28 else "000000000000" when X = 13 AND Y = 28 else "000000000000" when X = 14 AND Y = 28 else "000100000010" when X = 15 AND Y = 28 else "011000001001" when X = 16 AND Y = 28 else "011100001001" when X = 17 AND Y = 28 else "011100001001" when X = 18 AND Y = 28 else "011100001001" when X = 19 AND Y = 28 else "011100001001" when X = 20 AND Y = 28 else "011100001001" when X = 21 AND Y = 28 else "011100001001" when X = 22 AND Y = 28 else "011100001001" when X = 23 AND Y = 28 else "011100001001" when X = 24 AND Y = 28 else "011100001001" when X = 25 AND Y = 28 else "011100001001" when X = 26 AND Y = 28 else "010101001001" when X = 27 AND Y = 28 else "001110011001" when X = 28 AND Y = 28 else "100110011001" when X = 29 AND Y = 28 else "100110011001" when X = 30 AND Y = 28 else "100110011001" when X = 31 AND Y = 28 else "100110011001" when X = 32 AND Y = 28 else "100110011001" when X = 33 AND Y = 28 else "100110011001" when X = 34 AND Y = 28 else "100110011001" when X = 35 AND Y = 28 else "100110011001" when X = 36 AND Y = 28 else "100110011001" when X = 37 AND Y = 28 else "010110011001" when X = 38 AND Y = 28 else "010001011001" when X = 39 AND Y = 28 else "011100001001" when X = 40 AND Y = 28 else "011100001001" when X = 41 AND Y = 28 else "011100001001" when X = 42 AND Y = 28 else "011100001001" when X = 43 AND Y = 28 else "011100001001" when X = 44 AND Y = 28 else "011100001001" when X = 45 AND Y = 28 else "011100001001" when X = 46 AND Y = 28 else "011100001001" when X = 47 AND Y = 28 else "011100001001" when X = 48 AND Y = 28 else "011100001001" when X = 49 AND Y = 28 else "011100001010" when X = 50 AND Y = 28 else "010100000111" when X = 51 AND Y = 28 else "000000000000" when X = 52 AND Y = 28 else "000000000000" when X = 53 AND Y = 28 else "000000000000" when X = 54 AND Y = 28 else "000000000000" when X = 55 AND Y = 28 else "000000000000" when X = 56 AND Y = 28 else "000000000000" when X = 57 AND Y = 28 else "000000000000" when X = 58 AND Y = 28 else "000000000000" when X = 59 AND Y = 28 else "000000000000" when X = 60 AND Y = 28 else "000000000000" when X = 61 AND Y = 28 else "000000000000" when X = 62 AND Y = 28 else "001000100010" when X = 63 AND Y = 28 else "011110001001" when X = 64 AND Y = 28 else "111111110000" when X = 65 AND Y = 28 else "111111110000" when X = 66 AND Y = 28 else "111111110000" when X = 67 AND Y = 28 else "111111110000" when X = 68 AND Y = 28 else "111111110000" when X = 0 AND Y = 29 else "111111110000" when X = 1 AND Y = 29 else "101010111100" when X = 2 AND Y = 29 else "010101010101" when X = 3 AND Y = 29 else "000000000000" when X = 4 AND Y = 29 else "000000000000" when X = 5 AND Y = 29 else "000000000000" when X = 6 AND Y = 29 else "000000000000" when X = 7 AND Y = 29 else "000000000000" when X = 8 AND Y = 29 else "000000000000" when X = 9 AND Y = 29 else "000000000000" when X = 10 AND Y = 29 else "000000000000" when X = 11 AND Y = 29 else "000000000000" when X = 12 AND Y = 29 else "000000000000" when X = 13 AND Y = 29 else "000000000000" when X = 14 AND Y = 29 else "000100000010" when X = 15 AND Y = 29 else "011000001001" when X = 16 AND Y = 29 else "011000001001" when X = 17 AND Y = 29 else "001100001100" when X = 18 AND Y = 29 else "010001001010" when X = 19 AND Y = 29 else "010001101001" when X = 20 AND Y = 29 else "010001011001" when X = 21 AND Y = 29 else "010001101001" when X = 22 AND Y = 29 else "010001011001" when X = 23 AND Y = 29 else "011000101001" when X = 24 AND Y = 29 else "011100001001" when X = 25 AND Y = 29 else "011100001001" when X = 26 AND Y = 29 else "010101001001" when X = 27 AND Y = 29 else "001110011001" when X = 28 AND Y = 29 else "100110011001" when X = 29 AND Y = 29 else "011010011001" when X = 30 AND Y = 29 else "010110011001" when X = 31 AND Y = 29 else "010110011001" when X = 32 AND Y = 29 else "010110011001" when X = 33 AND Y = 29 else "010110011001" when X = 34 AND Y = 29 else "010110011001" when X = 35 AND Y = 29 else "010110011001" when X = 36 AND Y = 29 else "100010011001" when X = 37 AND Y = 29 else "010110011001" when X = 38 AND Y = 29 else "010001011001" when X = 39 AND Y = 29 else "011100001001" when X = 40 AND Y = 29 else "011100001001" when X = 41 AND Y = 29 else "011100001001" when X = 42 AND Y = 29 else "010101001001" when X = 43 AND Y = 29 else "010001101001" when X = 44 AND Y = 29 else "010001011001" when X = 45 AND Y = 29 else "010001011001" when X = 46 AND Y = 29 else "010001011001" when X = 47 AND Y = 29 else "001100101100" when X = 48 AND Y = 29 else "010100001011" when X = 49 AND Y = 29 else "011100001001" when X = 50 AND Y = 29 else "010100000111" when X = 51 AND Y = 29 else "000000000000" when X = 52 AND Y = 29 else "000000000000" when X = 53 AND Y = 29 else "000000000000" when X = 54 AND Y = 29 else "000000000000" when X = 55 AND Y = 29 else "000000000000" when X = 56 AND Y = 29 else "000000000000" when X = 57 AND Y = 29 else "000000000000" when X = 58 AND Y = 29 else "000000000000" when X = 59 AND Y = 29 else "000000000000" when X = 60 AND Y = 29 else "000000000000" when X = 61 AND Y = 29 else "000000000000" when X = 62 AND Y = 29 else "001100110011" when X = 63 AND Y = 29 else "100110101011" when X = 64 AND Y = 29 else "111111110000" when X = 65 AND Y = 29 else "111111110000" when X = 66 AND Y = 29 else "111111110000" when X = 67 AND Y = 29 else "111111110000" when X = 68 AND Y = 29 else "111111110000" when X = 0 AND Y = 30 else "111111110000" when X = 1 AND Y = 30 else "101010111100" when X = 2 AND Y = 30 else "010101010101" when X = 3 AND Y = 30 else "000000000000" when X = 4 AND Y = 30 else "000000000000" when X = 5 AND Y = 30 else "000000000000" when X = 6 AND Y = 30 else "000000000000" when X = 7 AND Y = 30 else "000000000000" when X = 8 AND Y = 30 else "000000000000" when X = 9 AND Y = 30 else "000000000000" when X = 10 AND Y = 30 else "000000000000" when X = 11 AND Y = 30 else "000000000000" when X = 12 AND Y = 30 else "000000000000" when X = 13 AND Y = 30 else "000000000000" when X = 14 AND Y = 30 else "001000000010" when X = 15 AND Y = 30 else "011000001001" when X = 16 AND Y = 30 else "010000011100" when X = 17 AND Y = 30 else "000100111101" when X = 18 AND Y = 30 else "000001111010" when X = 19 AND Y = 30 else "000010011000" when X = 20 AND Y = 30 else "000010011000" when X = 21 AND Y = 30 else "000010011000" when X = 22 AND Y = 30 else "000110001000" when X = 23 AND Y = 30 else "011000101001" when X = 24 AND Y = 30 else "011100001001" when X = 25 AND Y = 30 else "011100001001" when X = 26 AND Y = 30 else "010101001001" when X = 27 AND Y = 30 else "001110011001" when X = 28 AND Y = 30 else "100010011001" when X = 29 AND Y = 30 else "001010011001" when X = 30 AND Y = 30 else "000010001000" when X = 31 AND Y = 30 else "000001111010" when X = 32 AND Y = 30 else "000001011011" when X = 33 AND Y = 30 else "000001101011" when X = 34 AND Y = 30 else "000010001001" when X = 35 AND Y = 30 else "000010001000" when X = 36 AND Y = 30 else "100010011001" when X = 37 AND Y = 30 else "010110011001" when X = 38 AND Y = 30 else "010001011001" when X = 39 AND Y = 30 else "011100001001" when X = 40 AND Y = 30 else "011100001001" when X = 41 AND Y = 30 else "011100001001" when X = 42 AND Y = 30 else "010001011001" when X = 43 AND Y = 30 else "000010011000" when X = 44 AND Y = 30 else "000010011000" when X = 45 AND Y = 30 else "000010011000" when X = 46 AND Y = 30 else "000010001001" when X = 47 AND Y = 30 else "000001011100" when X = 48 AND Y = 30 else "001100101100" when X = 49 AND Y = 30 else "010100001011" when X = 50 AND Y = 30 else "010100000110" when X = 51 AND Y = 30 else "000000000000" when X = 52 AND Y = 30 else "000000000000" when X = 53 AND Y = 30 else "000000000000" when X = 54 AND Y = 30 else "000000000000" when X = 55 AND Y = 30 else "000000000000" when X = 56 AND Y = 30 else "000000000000" when X = 57 AND Y = 30 else "000000000000" when X = 58 AND Y = 30 else "000000000000" when X = 59 AND Y = 30 else "000000000000" when X = 60 AND Y = 30 else "000000000000" when X = 61 AND Y = 30 else "000000000000" when X = 62 AND Y = 30 else "001100110011" when X = 63 AND Y = 30 else "100110101011" when X = 64 AND Y = 30 else "111111110000" when X = 65 AND Y = 30 else "111111110000" when X = 66 AND Y = 30 else "111111110000" when X = 67 AND Y = 30 else "111111110000" when X = 68 AND Y = 30 else "111111110000" when X = 0 AND Y = 31 else "111111110000" when X = 1 AND Y = 31 else "100010101010" when X = 2 AND Y = 31 else "010001000100" when X = 3 AND Y = 31 else "000000000000" when X = 4 AND Y = 31 else "000000000000" when X = 5 AND Y = 31 else "000000000000" when X = 6 AND Y = 31 else "000000000000" when X = 7 AND Y = 31 else "000000000000" when X = 8 AND Y = 31 else "000000000000" when X = 9 AND Y = 31 else "000000000000" when X = 10 AND Y = 31 else "000000000000" when X = 11 AND Y = 31 else "000000000000" when X = 12 AND Y = 31 else "000000000000" when X = 13 AND Y = 31 else "000000000000" when X = 14 AND Y = 31 else "000100000011" when X = 15 AND Y = 31 else "010000001011" when X = 16 AND Y = 31 else "000100011111" when X = 17 AND Y = 31 else "000001111010" when X = 18 AND Y = 31 else "000010011000" when X = 19 AND Y = 31 else "000010001000" when X = 20 AND Y = 31 else "000010011000" when X = 21 AND Y = 31 else "000010001001" when X = 22 AND Y = 31 else "000101101010" when X = 23 AND Y = 31 else "010000101011" when X = 24 AND Y = 31 else "010100001011" when X = 25 AND Y = 31 else "011000001010" when X = 26 AND Y = 31 else "010101001001" when X = 27 AND Y = 31 else "001110011001" when X = 28 AND Y = 31 else "100010011001" when X = 29 AND Y = 31 else "001010011001" when X = 30 AND Y = 31 else "000010011000" when X = 31 AND Y = 31 else "000001001101" when X = 32 AND Y = 31 else "000100001111" when X = 33 AND Y = 31 else "000000111110" when X = 34 AND Y = 31 else "000010001001" when X = 35 AND Y = 31 else "000110011000" when X = 36 AND Y = 31 else "100010011001" when X = 37 AND Y = 31 else "010110011001" when X = 38 AND Y = 31 else "010001011001" when X = 39 AND Y = 31 else "011000001001" when X = 40 AND Y = 31 else "010100001011" when X = 41 AND Y = 31 else "010100001011" when X = 42 AND Y = 31 else "001101001011" when X = 43 AND Y = 31 else "000010001010" when X = 44 AND Y = 31 else "000010011000" when X = 45 AND Y = 31 else "000010001000" when X = 46 AND Y = 31 else "000010001000" when X = 47 AND Y = 31 else "000010011000" when X = 48 AND Y = 31 else "000001001101" when X = 49 AND Y = 31 else "001000001110" when X = 50 AND Y = 31 else "001100001000" when X = 51 AND Y = 31 else "000000000000" when X = 52 AND Y = 31 else "000000000000" when X = 53 AND Y = 31 else "000000000000" when X = 54 AND Y = 31 else "000000000000" when X = 55 AND Y = 31 else "000000000000" when X = 56 AND Y = 31 else "000000000000" when X = 57 AND Y = 31 else "000000000000" when X = 58 AND Y = 31 else "000000000000" when X = 59 AND Y = 31 else "000000000000" when X = 60 AND Y = 31 else "000000000000" when X = 61 AND Y = 31 else "000000000000" when X = 62 AND Y = 31 else "001000100010" when X = 63 AND Y = 31 else "011110001001" when X = 64 AND Y = 31 else "111111110000" when X = 65 AND Y = 31 else "111111110000" when X = 66 AND Y = 31 else "111111110000" when X = 67 AND Y = 31 else "111111110000" when X = 68 AND Y = 31 else "111111110000" when X = 0 AND Y = 32 else "111111110000" when X = 1 AND Y = 32 else "001101010101" when X = 2 AND Y = 32 else "000000000000" when X = 3 AND Y = 32 else "000000000000" when X = 4 AND Y = 32 else "000000000000" when X = 5 AND Y = 32 else "000000000000" when X = 6 AND Y = 32 else "000000000000" when X = 7 AND Y = 32 else "000000000000" when X = 8 AND Y = 32 else "000000000000" when X = 9 AND Y = 32 else "000000000000" when X = 10 AND Y = 32 else "000000000000" when X = 11 AND Y = 32 else "000000000000" when X = 12 AND Y = 32 else "000000000000" when X = 13 AND Y = 32 else "000000000000" when X = 14 AND Y = 32 else "000000000100" when X = 15 AND Y = 32 else "000100101111" when X = 16 AND Y = 32 else "000100011111" when X = 17 AND Y = 32 else "000001101011" when X = 18 AND Y = 32 else "000010001001" when X = 19 AND Y = 32 else "000010011000" when X = 20 AND Y = 32 else "000010001001" when X = 21 AND Y = 32 else "000001111010" when X = 22 AND Y = 32 else "000100011111" when X = 23 AND Y = 32 else "000100001111" when X = 24 AND Y = 32 else "000100001111" when X = 25 AND Y = 32 else "001100001101" when X = 26 AND Y = 32 else "010101001001" when X = 27 AND Y = 32 else "001110011001" when X = 28 AND Y = 32 else "100010011001" when X = 29 AND Y = 32 else "001010011001" when X = 30 AND Y = 32 else "000010011000" when X = 31 AND Y = 32 else "000001011100" when X = 32 AND Y = 32 else "000100011111" when X = 33 AND Y = 32 else "000001001101" when X = 34 AND Y = 32 else "000010001001" when X = 35 AND Y = 32 else "000110011000" when X = 36 AND Y = 32 else "100010011001" when X = 37 AND Y = 32 else "010110011001" when X = 38 AND Y = 32 else "010001011001" when X = 39 AND Y = 32 else "010100001011" when X = 40 AND Y = 32 else "000100001111" when X = 41 AND Y = 32 else "000100001111" when X = 42 AND Y = 32 else "000100001111" when X = 43 AND Y = 32 else "000001001101" when X = 44 AND Y = 32 else "000010001001" when X = 45 AND Y = 32 else "000010001000" when X = 46 AND Y = 32 else "000010001000" when X = 47 AND Y = 32 else "000010001001" when X = 48 AND Y = 32 else "000001001101" when X = 49 AND Y = 32 else "000100011111" when X = 50 AND Y = 32 else "000100011011" when X = 51 AND Y = 32 else "000000000000" when X = 52 AND Y = 32 else "000000000000" when X = 53 AND Y = 32 else "000000000000" when X = 54 AND Y = 32 else "000000000000" when X = 55 AND Y = 32 else "000000000000" when X = 56 AND Y = 32 else "000000000000" when X = 57 AND Y = 32 else "000000000000" when X = 58 AND Y = 32 else "000000000000" when X = 59 AND Y = 32 else "000000000000" when X = 60 AND Y = 32 else "000000000000" when X = 61 AND Y = 32 else "000000000000" when X = 62 AND Y = 32 else "000000000000" when X = 63 AND Y = 32 else "001000110011" when X = 64 AND Y = 32 else "111111110000" when X = 65 AND Y = 32 else "111111110000" when X = 66 AND Y = 32 else "111111110000" when X = 67 AND Y = 32 else "111111110000" when X = 68 AND Y = 32 else "111111110000" when X = 0 AND Y = 33 else "111111110000" when X = 1 AND Y = 33 else "001101010101" when X = 2 AND Y = 33 else "000000000000" when X = 3 AND Y = 33 else "000000000000" when X = 4 AND Y = 33 else "000000000000" when X = 5 AND Y = 33 else "000000000000" when X = 6 AND Y = 33 else "000000000000" when X = 7 AND Y = 33 else "000000000000" when X = 8 AND Y = 33 else "000000000000" when X = 9 AND Y = 33 else "000000000000" when X = 10 AND Y = 33 else "000000000000" when X = 11 AND Y = 33 else "000000000000" when X = 12 AND Y = 33 else "000000000000" when X = 13 AND Y = 33 else "000000000000" when X = 14 AND Y = 33 else "001000110100" when X = 15 AND Y = 33 else "011110101110" when X = 16 AND Y = 33 else "000100101111" when X = 17 AND Y = 33 else "000100011111" when X = 18 AND Y = 33 else "000001101011" when X = 19 AND Y = 33 else "000010011000" when X = 20 AND Y = 33 else "000001101010" when X = 21 AND Y = 33 else "000100011111" when X = 22 AND Y = 33 else "000100001111" when X = 23 AND Y = 33 else "000100001111" when X = 24 AND Y = 33 else "000100001111" when X = 25 AND Y = 33 else "000100001111" when X = 26 AND Y = 33 else "000101001101" when X = 27 AND Y = 33 else "001110011001" when X = 28 AND Y = 33 else "100010011001" when X = 29 AND Y = 33 else "001010011001" when X = 30 AND Y = 33 else "000010001000" when X = 31 AND Y = 33 else "000010001001" when X = 32 AND Y = 33 else "000010001001" when X = 33 AND Y = 33 else "000010001001" when X = 34 AND Y = 33 else "000010001000" when X = 35 AND Y = 33 else "000110011001" when X = 36 AND Y = 33 else "100010011001" when X = 37 AND Y = 33 else "010110011001" when X = 38 AND Y = 33 else "000001011011" when X = 39 AND Y = 33 else "000100001111" when X = 40 AND Y = 33 else "000100001111" when X = 41 AND Y = 33 else "000100001111" when X = 42 AND Y = 33 else "000100001111" when X = 43 AND Y = 33 else "000100001111" when X = 44 AND Y = 33 else "000001001101" when X = 45 AND Y = 33 else "000010001001" when X = 46 AND Y = 33 else "000010001001" when X = 47 AND Y = 33 else "000000111101" when X = 48 AND Y = 33 else "000100001111" when X = 49 AND Y = 33 else "001101101111" when X = 50 AND Y = 33 else "011010001010" when X = 51 AND Y = 33 else "000000000000" when X = 52 AND Y = 33 else "000000000000" when X = 53 AND Y = 33 else "000000000000" when X = 54 AND Y = 33 else "000000000000" when X = 55 AND Y = 33 else "000000000000" when X = 56 AND Y = 33 else "000000000000" when X = 57 AND Y = 33 else "000000000000" when X = 58 AND Y = 33 else "000000000000" when X = 59 AND Y = 33 else "000000000000" when X = 60 AND Y = 33 else "000000000000" when X = 61 AND Y = 33 else "000000000000" when X = 62 AND Y = 33 else "000000000000" when X = 63 AND Y = 33 else "001000100011" when X = 64 AND Y = 33 else "111111110000" when X = 65 AND Y = 33 else "111111110000" when X = 66 AND Y = 33 else "111111110000" when X = 67 AND Y = 33 else "111111110000" when X = 68 AND Y = 33 else "111111110000" when X = 0 AND Y = 34 else "111111110000" when X = 1 AND Y = 34 else "001101010101" when X = 2 AND Y = 34 else "000000000000" when X = 3 AND Y = 34 else "000000000000" when X = 4 AND Y = 34 else "000000000000" when X = 5 AND Y = 34 else "000000000000" when X = 6 AND Y = 34 else "000000000000" when X = 7 AND Y = 34 else "000000000000" when X = 8 AND Y = 34 else "000000000000" when X = 9 AND Y = 34 else "000000000000" when X = 10 AND Y = 34 else "000000000000" when X = 11 AND Y = 34 else "000000000000" when X = 12 AND Y = 34 else "000000000000" when X = 13 AND Y = 34 else "000000000000" when X = 14 AND Y = 34 else "001000110100" when X = 15 AND Y = 34 else "111111110000" when X = 16 AND Y = 34 else "011110101111" when X = 17 AND Y = 34 else "000100111111" when X = 18 AND Y = 34 else "000100101111" when X = 19 AND Y = 34 else "000001101011" when X = 20 AND Y = 34 else "000001101011" when X = 21 AND Y = 34 else "000100001111" when X = 22 AND Y = 34 else "000100001111" when X = 23 AND Y = 34 else "000100001111" when X = 24 AND Y = 34 else "000100001111" when X = 25 AND Y = 34 else "000100001111" when X = 26 AND Y = 34 else "000001001101" when X = 27 AND Y = 34 else "001110011001" when X = 28 AND Y = 34 else "100010011001" when X = 29 AND Y = 34 else "001010011001" when X = 30 AND Y = 34 else "000010001000" when X = 31 AND Y = 34 else "000010001000" when X = 32 AND Y = 34 else "000010011000" when X = 33 AND Y = 34 else "000010001000" when X = 34 AND Y = 34 else "000010001000" when X = 35 AND Y = 34 else "000010011000" when X = 36 AND Y = 34 else "100010011001" when X = 37 AND Y = 34 else "010110011001" when X = 38 AND Y = 34 else "000001011100" when X = 39 AND Y = 34 else "000100001111" when X = 40 AND Y = 34 else "000100001111" when X = 41 AND Y = 34 else "000100001111" when X = 42 AND Y = 34 else "000100001111" when X = 43 AND Y = 34 else "000100001111" when X = 44 AND Y = 34 else "000000111110" when X = 45 AND Y = 34 else "000010001001" when X = 46 AND Y = 34 else "000000111101" when X = 47 AND Y = 34 else "000100001111" when X = 48 AND Y = 34 else "010001111111" when X = 49 AND Y = 34 else "101011011101" when X = 50 AND Y = 34 else "011010011010" when X = 51 AND Y = 34 else "000000000000" when X = 52 AND Y = 34 else "000000000000" when X = 53 AND Y = 34 else "000000000000" when X = 54 AND Y = 34 else "000000000000" when X = 55 AND Y = 34 else "000000000000" when X = 56 AND Y = 34 else "000000000000" when X = 57 AND Y = 34 else "000000000000" when X = 58 AND Y = 34 else "000000000000" when X = 59 AND Y = 34 else "000000000000" when X = 60 AND Y = 34 else "000000000000" when X = 61 AND Y = 34 else "000000000000" when X = 62 AND Y = 34 else "000000000000" when X = 63 AND Y = 34 else "001000100011" when X = 64 AND Y = 34 else "111111110000" when X = 65 AND Y = 34 else "111111110000" when X = 66 AND Y = 34 else "111111110000" when X = 67 AND Y = 34 else "111111110000" when X = 68 AND Y = 34 else "111111110000" when X = 0 AND Y = 35 else "111111110000" when X = 1 AND Y = 35 else "001101010101" when X = 2 AND Y = 35 else "000000000000" when X = 3 AND Y = 35 else "000000000000" when X = 4 AND Y = 35 else "000000000000" when X = 5 AND Y = 35 else "000000000000" when X = 6 AND Y = 35 else "000000000000" when X = 7 AND Y = 35 else "000000000000" when X = 8 AND Y = 35 else "000000000000" when X = 9 AND Y = 35 else "000000000000" when X = 10 AND Y = 35 else "000000000000" when X = 11 AND Y = 35 else "000000000000" when X = 12 AND Y = 35 else "000000000000" when X = 13 AND Y = 35 else "000000000000" when X = 14 AND Y = 35 else "001000110100" when X = 15 AND Y = 35 else "111111110000" when X = 16 AND Y = 35 else "111111110000" when X = 17 AND Y = 35 else "011010011111" when X = 18 AND Y = 35 else "001000111111" when X = 19 AND Y = 35 else "000100101110" when X = 20 AND Y = 35 else "000000111110" when X = 21 AND Y = 35 else "000100001111" when X = 22 AND Y = 35 else "000100001111" when X = 23 AND Y = 35 else "000100001111" when X = 24 AND Y = 35 else "000100001111" when X = 25 AND Y = 35 else "000100001111" when X = 26 AND Y = 35 else "000001001101" when X = 27 AND Y = 35 else "001110011001" when X = 28 AND Y = 35 else "100110011001" when X = 29 AND Y = 35 else "011110011001" when X = 30 AND Y = 35 else "011010011001" when X = 31 AND Y = 35 else "011010011001" when X = 32 AND Y = 35 else "011010011001" when X = 33 AND Y = 35 else "011010011001" when X = 34 AND Y = 35 else "011010011001" when X = 35 AND Y = 35 else "011010011001" when X = 36 AND Y = 35 else "100110011001" when X = 37 AND Y = 35 else "010110011001" when X = 38 AND Y = 35 else "000001011100" when X = 39 AND Y = 35 else "000100001111" when X = 40 AND Y = 35 else "000100001111" when X = 41 AND Y = 35 else "000100001111" when X = 42 AND Y = 35 else "000100001111" when X = 43 AND Y = 35 else "000100001111" when X = 44 AND Y = 35 else "000100011111" when X = 45 AND Y = 35 else "000000111101" when X = 46 AND Y = 35 else "000100001111" when X = 47 AND Y = 35 else "010001101111" when X = 48 AND Y = 35 else "100011001110" when X = 49 AND Y = 35 else "111111110000" when X = 50 AND Y = 35 else "011010011010" when X = 51 AND Y = 35 else "000000000000" when X = 52 AND Y = 35 else "000000000000" when X = 53 AND Y = 35 else "000000000000" when X = 54 AND Y = 35 else "000000000000" when X = 55 AND Y = 35 else "000000000000" when X = 56 AND Y = 35 else "000000000000" when X = 57 AND Y = 35 else "000000000000" when X = 58 AND Y = 35 else "000000000000" when X = 59 AND Y = 35 else "000000000000" when X = 60 AND Y = 35 else "000000000000" when X = 61 AND Y = 35 else "000000000000" when X = 62 AND Y = 35 else "000000000000" when X = 63 AND Y = 35 else "001000100011" when X = 64 AND Y = 35 else "111111110000" when X = 65 AND Y = 35 else "111111110000" when X = 66 AND Y = 35 else "111111110000" when X = 67 AND Y = 35 else "111111110000" when X = 68 AND Y = 35 else "111111110000" when X = 0 AND Y = 36 else "111111110000" when X = 1 AND Y = 36 else "001101010101" when X = 2 AND Y = 36 else "000000000000" when X = 3 AND Y = 36 else "000000000000" when X = 4 AND Y = 36 else "000000000000" when X = 5 AND Y = 36 else "000000000000" when X = 6 AND Y = 36 else "000000000000" when X = 7 AND Y = 36 else "000000000000" when X = 8 AND Y = 36 else "000000000000" when X = 9 AND Y = 36 else "000000000000" when X = 10 AND Y = 36 else "000000000000" when X = 11 AND Y = 36 else "000000000000" when X = 12 AND Y = 36 else "000000000000" when X = 13 AND Y = 36 else "000000000000" when X = 14 AND Y = 36 else "001000110100" when X = 15 AND Y = 36 else "111111110000" when X = 16 AND Y = 36 else "111111110000" when X = 17 AND Y = 36 else "111111110000" when X = 18 AND Y = 36 else "010110011111" when X = 19 AND Y = 36 else "001101101111" when X = 20 AND Y = 36 else "001101101111" when X = 21 AND Y = 36 else "001101011111" when X = 22 AND Y = 36 else "000100001111" when X = 23 AND Y = 36 else "000100001111" when X = 24 AND Y = 36 else "000100001111" when X = 25 AND Y = 36 else "001000111111" when X = 26 AND Y = 36 else "010010001110" when X = 27 AND Y = 36 else "011010111011" when X = 28 AND Y = 36 else "100110111011" when X = 29 AND Y = 36 else "100110111011" when X = 30 AND Y = 36 else "100110111011" when X = 31 AND Y = 36 else "100110111011" when X = 32 AND Y = 36 else "100110111011" when X = 33 AND Y = 36 else "100110111011" when X = 34 AND Y = 36 else "100110111011" when X = 35 AND Y = 36 else "100110111011" when X = 36 AND Y = 36 else "100110111011" when X = 37 AND Y = 36 else "011010111011" when X = 38 AND Y = 36 else "010010001101" when X = 39 AND Y = 36 else "001101101111" when X = 40 AND Y = 36 else "000100011111" when X = 41 AND Y = 36 else "000100001111" when X = 42 AND Y = 36 else "000100001111" when X = 43 AND Y = 36 else "000100111111" when X = 44 AND Y = 36 else "001101101111" when X = 45 AND Y = 36 else "001101101111" when X = 46 AND Y = 36 else "010001101111" when X = 47 AND Y = 36 else "100011001110" when X = 48 AND Y = 36 else "111111110000" when X = 49 AND Y = 36 else "111111110000" when X = 50 AND Y = 36 else "011010011010" when X = 51 AND Y = 36 else "000000000000" when X = 52 AND Y = 36 else "000000000000" when X = 53 AND Y = 36 else "000000000000" when X = 54 AND Y = 36 else "000000000000" when X = 55 AND Y = 36 else "000000000000" when X = 56 AND Y = 36 else "000000000000" when X = 57 AND Y = 36 else "000000000000" when X = 58 AND Y = 36 else "000000000000" when X = 59 AND Y = 36 else "000000000000" when X = 60 AND Y = 36 else "000000000000" when X = 61 AND Y = 36 else "000000000000" when X = 62 AND Y = 36 else "000000000000" when X = 63 AND Y = 36 else "001000100011" when X = 64 AND Y = 36 else "111111110000" when X = 65 AND Y = 36 else "111111110000" when X = 66 AND Y = 36 else "111111110000" when X = 67 AND Y = 36 else "111111110000" when X = 68 AND Y = 36 else "111111110000" when X = 0 AND Y = 37 else "111111110000" when X = 1 AND Y = 37 else "010101111000" when X = 2 AND Y = 37 else "000100010001" when X = 3 AND Y = 37 else "000000000000" when X = 4 AND Y = 37 else "000000000000" when X = 5 AND Y = 37 else "000000000000" when X = 6 AND Y = 37 else "000000000000" when X = 7 AND Y = 37 else "000000000000" when X = 8 AND Y = 37 else "000000000000" when X = 9 AND Y = 37 else "000000000000" when X = 10 AND Y = 37 else "000000000000" when X = 11 AND Y = 37 else "000000000000" when X = 12 AND Y = 37 else "000000000000" when X = 13 AND Y = 37 else "000000010001" when X = 14 AND Y = 37 else "010001100110" when X = 15 AND Y = 37 else "111111110000" when X = 16 AND Y = 37 else "111111110000" when X = 17 AND Y = 37 else "111111110000" when X = 18 AND Y = 37 else "111111110000" when X = 19 AND Y = 37 else "111111110000" when X = 20 AND Y = 37 else "111111110000" when X = 21 AND Y = 37 else "100011001110" when X = 22 AND Y = 37 else "001001011111" when X = 23 AND Y = 37 else "001001001111" when X = 24 AND Y = 37 else "001001001111" when X = 25 AND Y = 37 else "011010011111" when X = 26 AND Y = 37 else "111111110000" when X = 27 AND Y = 37 else "111111110000" when X = 28 AND Y = 37 else "111111110000" when X = 29 AND Y = 37 else "111111110000" when X = 30 AND Y = 37 else "111111110000" when X = 31 AND Y = 37 else "111111110000" when X = 32 AND Y = 37 else "111111110000" when X = 33 AND Y = 37 else "111111110000" when X = 34 AND Y = 37 else "111111110000" when X = 35 AND Y = 37 else "111111110000" when X = 36 AND Y = 37 else "111111110000" when X = 37 AND Y = 37 else "111111110000" when X = 38 AND Y = 37 else "111111110000" when X = 39 AND Y = 37 else "111111110000" when X = 40 AND Y = 37 else "001101011111" when X = 41 AND Y = 37 else "001001001111" when X = 42 AND Y = 37 else "001001001111" when X = 43 AND Y = 37 else "010110001111" when X = 44 AND Y = 37 else "111111110000" when X = 45 AND Y = 37 else "111111110000" when X = 46 AND Y = 37 else "111111110000" when X = 47 AND Y = 37 else "111111110000" when X = 48 AND Y = 37 else "111111110000" when X = 49 AND Y = 37 else "111111110000" when X = 50 AND Y = 37 else "011110101011" when X = 51 AND Y = 37 else "001000110011" when X = 52 AND Y = 37 else "000000000000" when X = 53 AND Y = 37 else "000000000000" when X = 54 AND Y = 37 else "000000000000" when X = 55 AND Y = 37 else "000000000000" when X = 56 AND Y = 37 else "000000000000" when X = 57 AND Y = 37 else "000000000000" when X = 58 AND Y = 37 else "000000000000" when X = 59 AND Y = 37 else "000000000000" when X = 60 AND Y = 37 else "000000000000" when X = 61 AND Y = 37 else "000000000000" when X = 62 AND Y = 37 else "000000010001" when X = 63 AND Y = 37 else "001101010110" when X = 64 AND Y = 37 else "111111110000" when X = 65 AND Y = 37 else "111111110000" when X = 66 AND Y = 37 else "111111110000" when X = 67 AND Y = 37 else "111111110000" when X = 68 AND Y = 37 else "111111110000" when X = 0 AND Y = 38 else "111111110000" when X = 1 AND Y = 38 else "111111110000" when X = 2 AND Y = 38 else "010110001000" when X = 3 AND Y = 38 else "000100010001" when X = 4 AND Y = 38 else "000100010001" when X = 5 AND Y = 38 else "000100010001" when X = 6 AND Y = 38 else "000100010001" when X = 7 AND Y = 38 else "000100010001" when X = 8 AND Y = 38 else "000100010001" when X = 9 AND Y = 38 else "000100010001" when X = 10 AND Y = 38 else "000100010001" when X = 11 AND Y = 38 else "000100010001" when X = 12 AND Y = 38 else "000100010001" when X = 13 AND Y = 38 else "010001100111" when X = 14 AND Y = 38 else "111111110000" when X = 15 AND Y = 38 else "111111110000" when X = 16 AND Y = 38 else "111111110000" when X = 17 AND Y = 38 else "111111110000" when X = 18 AND Y = 38 else "111111110000" when X = 19 AND Y = 38 else "111111110000" when X = 20 AND Y = 38 else "111111110000" when X = 21 AND Y = 38 else "111111110000" when X = 22 AND Y = 38 else "111111110000" when X = 23 AND Y = 38 else "111111110000" when X = 24 AND Y = 38 else "111111110000" when X = 25 AND Y = 38 else "111111110000" when X = 26 AND Y = 38 else "111111110000" when X = 27 AND Y = 38 else "111111110000" when X = 28 AND Y = 38 else "111111110000" when X = 29 AND Y = 38 else "111111110000" when X = 30 AND Y = 38 else "111111110000" when X = 31 AND Y = 38 else "111111110000" when X = 32 AND Y = 38 else "111111110000" when X = 33 AND Y = 38 else "111111110000" when X = 34 AND Y = 38 else "111111110000" when X = 35 AND Y = 38 else "111111110000" when X = 36 AND Y = 38 else "111111110000" when X = 37 AND Y = 38 else "111111110000" when X = 38 AND Y = 38 else "111111110000" when X = 39 AND Y = 38 else "111111110000" when X = 40 AND Y = 38 else "111111110000" when X = 41 AND Y = 38 else "111111110000" when X = 42 AND Y = 38 else "111111110000" when X = 43 AND Y = 38 else "111111110000" when X = 44 AND Y = 38 else "111111110000" when X = 45 AND Y = 38 else "111111110000" when X = 46 AND Y = 38 else "111111110000" when X = 47 AND Y = 38 else "111111110000" when X = 48 AND Y = 38 else "111111110000" when X = 49 AND Y = 38 else "111111110000" when X = 50 AND Y = 38 else "111111110000" when X = 51 AND Y = 38 else "100010111100" when X = 52 AND Y = 38 else "000100100010" when X = 53 AND Y = 38 else "000100010001" when X = 54 AND Y = 38 else "000100010001" when X = 55 AND Y = 38 else "000100010001" when X = 56 AND Y = 38 else "000100010001" when X = 57 AND Y = 38 else "000100010001" when X = 58 AND Y = 38 else "000100010001" when X = 59 AND Y = 38 else "000100010001" when X = 60 AND Y = 38 else "000100010001" when X = 61 AND Y = 38 else "000100010001" when X = 62 AND Y = 38 else "010001010110" when X = 63 AND Y = 38 else "111111110000" when X = 64 AND Y = 38 else "111111110000" when X = 65 AND Y = 38 else "111111110000" when X = 66 AND Y = 38 else "111111110000" when X = 67 AND Y = 38 else "111111110000" when X = 68 AND Y = 38 else "111111110000" when X = 0 AND Y = 39 else "111111110000" when X = 1 AND Y = 39 else "111111110000" when X = 2 AND Y = 39 else "111111110101" when X = 3 AND Y = 39 else "100011001100" when X = 4 AND Y = 39 else "100011001100" when X = 5 AND Y = 39 else "100011001100" when X = 6 AND Y = 39 else "100011001100" when X = 7 AND Y = 39 else "100011001100" when X = 8 AND Y = 39 else "100011001100" when X = 9 AND Y = 39 else "100011001100" when X = 10 AND Y = 39 else "100011001100" when X = 11 AND Y = 39 else "100011001100" when X = 12 AND Y = 39 else "100010111100" when X = 13 AND Y = 39 else "110011101010" when X = 14 AND Y = 39 else "111111110000" when X = 15 AND Y = 39 else "111111110000" when X = 16 AND Y = 39 else "111111110000" when X = 17 AND Y = 39 else "111111110000" when X = 18 AND Y = 39 else "111111110000" when X = 19 AND Y = 39 else "111111110000" when X = 20 AND Y = 39 else "111111110000" when X = 21 AND Y = 39 else "111111110000" when X = 22 AND Y = 39 else "111111110000" when X = 23 AND Y = 39 else "111111110000" when X = 24 AND Y = 39 else "111111110000" when X = 25 AND Y = 39 else "111111110000" when X = 26 AND Y = 39 else "111111110000" when X = 27 AND Y = 39 else "111111110000" when X = 28 AND Y = 39 else "111111110000" when X = 29 AND Y = 39 else "111111110000" when X = 30 AND Y = 39 else "111111110000" when X = 31 AND Y = 39 else "111111110000" when X = 32 AND Y = 39 else "111111110000" when X = 33 AND Y = 39 else "111111110000" when X = 34 AND Y = 39 else "111111110000" when X = 35 AND Y = 39 else "111111110000" when X = 36 AND Y = 39 else "111111110000" when X = 37 AND Y = 39 else "111111110000" when X = 38 AND Y = 39 else "111111110000" when X = 39 AND Y = 39 else "111111110000" when X = 40 AND Y = 39 else "111111110000" when X = 41 AND Y = 39 else "111111110000" when X = 42 AND Y = 39 else "111111110000" when X = 43 AND Y = 39 else "111111110000" when X = 44 AND Y = 39 else "111111110000" when X = 45 AND Y = 39 else "111111110000" when X = 46 AND Y = 39 else "111111110000" when X = 47 AND Y = 39 else "111111110000" when X = 48 AND Y = 39 else "111111110000" when X = 49 AND Y = 39 else "111111110000" when X = 50 AND Y = 39 else "111111110000" when X = 51 AND Y = 39 else "111111110000" when X = 52 AND Y = 39 else "100011001101" when X = 53 AND Y = 39 else "100011001100" when X = 54 AND Y = 39 else "100011001100" when X = 55 AND Y = 39 else "100011001100" when X = 56 AND Y = 39 else "100011001100" when X = 57 AND Y = 39 else "100011001100" when X = 58 AND Y = 39 else "100011001100" when X = 59 AND Y = 39 else "100011001100" when X = 60 AND Y = 39 else "100011001100" when X = 61 AND Y = 39 else "100010111100" when X = 62 AND Y = 39 else "101011011100" when X = 63 AND Y = 39 else "111111110000" when X = 64 AND Y = 39 else "111111110000" when X = 65 AND Y = 39 else "111111110000" when X = 66 AND Y = 39 else "111111110000" when X = 67 AND Y = 39 else "111111110000" when X = 68 AND Y = 39 else "111111110000" when X = 0 AND Y = 40 else "111111110000" when X = 1 AND Y = 40 else "111111110000" when X = 2 AND Y = 40 else "111111110000" when X = 3 AND Y = 40 else "111111110000" when X = 4 AND Y = 40 else "111111110000" when X = 5 AND Y = 40 else "111111110000" when X = 6 AND Y = 40 else "111111110000" when X = 7 AND Y = 40 else "111111110000" when X = 8 AND Y = 40 else "111111110000" when X = 9 AND Y = 40 else "111111110000" when X = 10 AND Y = 40 else "111111110000" when X = 11 AND Y = 40 else "111111110000" when X = 12 AND Y = 40 else "111111110000" when X = 13 AND Y = 40 else "111111110000" when X = 14 AND Y = 40 else "111111110000" when X = 15 AND Y = 40 else "111111110000" when X = 16 AND Y = 40 else "111111110000" when X = 17 AND Y = 40 else "111111110000" when X = 18 AND Y = 40 else "111111110000" when X = 19 AND Y = 40 else "111111110000" when X = 20 AND Y = 40 else "111111110000" when X = 21 AND Y = 40 else "111111110000" when X = 22 AND Y = 40 else "111111110000" when X = 23 AND Y = 40 else "111111110000" when X = 24 AND Y = 40 else "111111110000" when X = 25 AND Y = 40 else "111111110000" when X = 26 AND Y = 40 else "111111110000" when X = 27 AND Y = 40 else "111111110000" when X = 28 AND Y = 40 else "111111110000" when X = 29 AND Y = 40 else "111111110000" when X = 30 AND Y = 40 else "111111110000" when X = 31 AND Y = 40 else "111111110000" when X = 32 AND Y = 40 else "111111110000" when X = 33 AND Y = 40 else "111111110000" when X = 34 AND Y = 40 else "111111110000" when X = 35 AND Y = 40 else "111111110000" when X = 36 AND Y = 40 else "111111110000" when X = 37 AND Y = 40 else "111111110000" when X = 38 AND Y = 40 else "111111110000" when X = 39 AND Y = 40 else "111111110000" when X = 40 AND Y = 40 else "111111110000" when X = 41 AND Y = 40 else "111111110000" when X = 42 AND Y = 40 else "111111110000" when X = 43 AND Y = 40 else "111111110000" when X = 44 AND Y = 40 else "111111110000" when X = 45 AND Y = 40 else "111111110000" when X = 46 AND Y = 40 else "111111110000" when X = 47 AND Y = 40 else "111111110000" when X = 48 AND Y = 40 else "111111110000" when X = 49 AND Y = 40 else "111111110000" when X = 50 AND Y = 40 else "111111110000" when X = 51 AND Y = 40 else "111111110000" when X = 52 AND Y = 40 else "111111110000" when X = 53 AND Y = 40 else "111111110000" when X = 54 AND Y = 40 else "111111110000" when X = 55 AND Y = 40 else "111111110000" when X = 56 AND Y = 40 else "111111110000" when X = 57 AND Y = 40 else "111111110000" when X = 58 AND Y = 40 else "111111110000" when X = 59 AND Y = 40 else "111111110000" when X = 60 AND Y = 40 else "111111110000" when X = 61 AND Y = 40 else "111111110000" when X = 62 AND Y = 40 else "111111110000" when X = 63 AND Y = 40 else "111111110000" when X = 64 AND Y = 40 else "111111110000" when X = 65 AND Y = 40 else "111111110000" when X = 66 AND Y = 40 else "111111110000" when X = 67 AND Y = 40 else "111111110000" when X = 68 AND Y = 40 else "111111110000" when X = 0 AND Y = 41 else "111111110000" when X = 1 AND Y = 41 else "111111110000" when X = 2 AND Y = 41 else "111111110000" when X = 3 AND Y = 41 else "111111110000" when X = 4 AND Y = 41 else "111111110000" when X = 5 AND Y = 41 else "111111110000" when X = 6 AND Y = 41 else "111111110000" when X = 7 AND Y = 41 else "111111110000" when X = 8 AND Y = 41 else "111111110000" when X = 9 AND Y = 41 else "111111110000" when X = 10 AND Y = 41 else "111111110000" when X = 11 AND Y = 41 else "111111110000" when X = 12 AND Y = 41 else "111111110000" when X = 13 AND Y = 41 else "111111110000" when X = 14 AND Y = 41 else "111111110000" when X = 15 AND Y = 41 else "111111110000" when X = 16 AND Y = 41 else "111111110000" when X = 17 AND Y = 41 else "111111110000" when X = 18 AND Y = 41 else "111111110000" when X = 19 AND Y = 41 else "111111110000" when X = 20 AND Y = 41 else "111111110000" when X = 21 AND Y = 41 else "111111110000" when X = 22 AND Y = 41 else "111111110000" when X = 23 AND Y = 41 else "111111110000" when X = 24 AND Y = 41 else "111111110000" when X = 25 AND Y = 41 else "111111110000" when X = 26 AND Y = 41 else "111111110000" when X = 27 AND Y = 41 else "111111110000" when X = 28 AND Y = 41 else "111111110000" when X = 29 AND Y = 41 else "111111110000" when X = 30 AND Y = 41 else "111111110000" when X = 31 AND Y = 41 else "111111110000" when X = 32 AND Y = 41 else "111111110000" when X = 33 AND Y = 41 else "111111110000" when X = 34 AND Y = 41 else "111111110000" when X = 35 AND Y = 41 else "111111110000" when X = 36 AND Y = 41 else "111111110000" when X = 37 AND Y = 41 else "111111110000" when X = 38 AND Y = 41 else "111111110000" when X = 39 AND Y = 41 else "111111110000" when X = 40 AND Y = 41 else "111111110000" when X = 41 AND Y = 41 else "111111110000" when X = 42 AND Y = 41 else "111111110000" when X = 43 AND Y = 41 else "111111110000" when X = 44 AND Y = 41 else "111111110000" when X = 45 AND Y = 41 else "111111110000" when X = 46 AND Y = 41 else "111111110000" when X = 47 AND Y = 41 else "111111110000" when X = 48 AND Y = 41 else "111111110000" when X = 49 AND Y = 41 else "111111110000" when X = 50 AND Y = 41 else "111111110000" when X = 51 AND Y = 41 else "111111110000" when X = 52 AND Y = 41 else "111111110000" when X = 53 AND Y = 41 else "111111110000" when X = 54 AND Y = 41 else "111111110000" when X = 55 AND Y = 41 else "111111110000" when X = 56 AND Y = 41 else "111111110000" when X = 57 AND Y = 41 else "111111110000" when X = 58 AND Y = 41 else "111111110000" when X = 59 AND Y = 41 else "111111110000" when X = 60 AND Y = 41 else "111111110000" when X = 61 AND Y = 41 else "111111110000" when X = 62 AND Y = 41 else "111111110000" when X = 63 AND Y = 41 else "111111110000" when X = 64 AND Y = 41 else "111111110000" when X = 65 AND Y = 41 else "111111110000" when X = 66 AND Y = 41 else "111111110000" when X = 67 AND Y = 41 else "111111110000" when X = 68 AND Y = 41 else "111111110000" when X = 0 AND Y = 42 else "111111110000" when X = 1 AND Y = 42 else "111111110000" when X = 2 AND Y = 42 else "111111110000" when X = 3 AND Y = 42 else "111111110000" when X = 4 AND Y = 42 else "111111110000" when X = 5 AND Y = 42 else "111111110000" when X = 6 AND Y = 42 else "111111110000" when X = 7 AND Y = 42 else "111111110000" when X = 8 AND Y = 42 else "111111110000" when X = 9 AND Y = 42 else "111111110000" when X = 10 AND Y = 42 else "111111110000" when X = 11 AND Y = 42 else "111111110000" when X = 12 AND Y = 42 else "111111110000" when X = 13 AND Y = 42 else "111111110000" when X = 14 AND Y = 42 else "111111110000" when X = 15 AND Y = 42 else "111111110000" when X = 16 AND Y = 42 else "111111110000" when X = 17 AND Y = 42 else "111111110000" when X = 18 AND Y = 42 else "111111110000" when X = 19 AND Y = 42 else "111111110000" when X = 20 AND Y = 42 else "111111110000" when X = 21 AND Y = 42 else "111111110000" when X = 22 AND Y = 42 else "111111110000" when X = 23 AND Y = 42 else "111111110000" when X = 24 AND Y = 42 else "111111110000" when X = 25 AND Y = 42 else "111111110000" when X = 26 AND Y = 42 else "111111110000" when X = 27 AND Y = 42 else "111111110000" when X = 28 AND Y = 42 else "111111110000" when X = 29 AND Y = 42 else "111111110000" when X = 30 AND Y = 42 else "111111110000" when X = 31 AND Y = 42 else "111111110000" when X = 32 AND Y = 42 else "111111110000" when X = 33 AND Y = 42 else "111111110000" when X = 34 AND Y = 42 else "111111110000" when X = 35 AND Y = 42 else "111111110000" when X = 36 AND Y = 42 else "111111110000" when X = 37 AND Y = 42 else "111111110000" when X = 38 AND Y = 42 else "111111110000" when X = 39 AND Y = 42 else "111111110000" when X = 40 AND Y = 42 else "111111110000" when X = 41 AND Y = 42 else "111111110000" when X = 42 AND Y = 42 else "111111110000" when X = 43 AND Y = 42 else "111111110000" when X = 44 AND Y = 42 else "111111110000" when X = 45 AND Y = 42 else "111111110000" when X = 46 AND Y = 42 else "111111110000" when X = 47 AND Y = 42 else "111111110000" when X = 48 AND Y = 42 else "111111110000" when X = 49 AND Y = 42 else "111111110000" when X = 50 AND Y = 42 else "111111110000" when X = 51 AND Y = 42 else "111111110000" when X = 52 AND Y = 42 else "111111110000" when X = 53 AND Y = 42 else "111111110000" when X = 54 AND Y = 42 else "111111110000" when X = 55 AND Y = 42 else "111111110000" when X = 56 AND Y = 42 else "111111110000" when X = 57 AND Y = 42 else "111111110000" when X = 58 AND Y = 42 else "111111110000" when X = 59 AND Y = 42 else "111111110000" when X = 60 AND Y = 42 else "111111110000" when X = 61 AND Y = 42 else "111111110000" when X = 62 AND Y = 42 else "111111110000" when X = 63 AND Y = 42 else "111111110000" when X = 64 AND Y = 42 else "111111110000" when X = 65 AND Y = 42 else "111111110000" when X = 66 AND Y = 42 else "111111110000" when X = 67 AND Y = 42 else "111111110000" when X = 68 AND Y = 42 else "111111110000" when X = 0 AND Y = 43 else "111111110000" when X = 1 AND Y = 43 else "111111110000" when X = 2 AND Y = 43 else "111111110000" when X = 3 AND Y = 43 else "111111110000" when X = 4 AND Y = 43 else "111111110000" when X = 5 AND Y = 43 else "111111110000" when X = 6 AND Y = 43 else "111111110000" when X = 7 AND Y = 43 else "111111110000" when X = 8 AND Y = 43 else "111111110000" when X = 9 AND Y = 43 else "111111110000" when X = 10 AND Y = 43 else "111111110000" when X = 11 AND Y = 43 else "111111110000" when X = 12 AND Y = 43 else "111111110000" when X = 13 AND Y = 43 else "111111110000" when X = 14 AND Y = 43 else "111111110000" when X = 15 AND Y = 43 else "111111110000" when X = 16 AND Y = 43 else "111111110000" when X = 17 AND Y = 43 else "111111110000" when X = 18 AND Y = 43 else "111111110000" when X = 19 AND Y = 43 else "111111110000" when X = 20 AND Y = 43 else "111111110000" when X = 21 AND Y = 43 else "111111110000" when X = 22 AND Y = 43 else "111111110000" when X = 23 AND Y = 43 else "111111110000" when X = 24 AND Y = 43 else "111111110000" when X = 25 AND Y = 43 else "111111110000" when X = 26 AND Y = 43 else "111111110000" when X = 27 AND Y = 43 else "111111110000" when X = 28 AND Y = 43 else "111111110000" when X = 29 AND Y = 43 else "111111110000" when X = 30 AND Y = 43 else "111111110000" when X = 31 AND Y = 43 else "111111110000" when X = 32 AND Y = 43 else "111111110000" when X = 33 AND Y = 43 else "111111110000" when X = 34 AND Y = 43 else "111111110000" when X = 35 AND Y = 43 else "111111110000" when X = 36 AND Y = 43 else "111111110000" when X = 37 AND Y = 43 else "111111110000" when X = 38 AND Y = 43 else "111111110000" when X = 39 AND Y = 43 else "111111110000" when X = 40 AND Y = 43 else "111111110000" when X = 41 AND Y = 43 else "111111110000" when X = 42 AND Y = 43 else "111111110000" when X = 43 AND Y = 43 else "111111110000" when X = 44 AND Y = 43 else "111111110000" when X = 45 AND Y = 43 else "111111110000" when X = 46 AND Y = 43 else "111111110000" when X = 47 AND Y = 43 else "111111110000" when X = 48 AND Y = 43 else "111111110000" when X = 49 AND Y = 43 else "111111110000" when X = 50 AND Y = 43 else "111111110000" when X = 51 AND Y = 43 else "111111110000" when X = 52 AND Y = 43 else "111111110000" when X = 53 AND Y = 43 else "111111110000" when X = 54 AND Y = 43 else "111111110000" when X = 55 AND Y = 43 else "111111110000" when X = 56 AND Y = 43 else "111111110000" when X = 57 AND Y = 43 else "111111110000" when X = 58 AND Y = 43 else "111111110000" when X = 59 AND Y = 43 else "111111110000" when X = 60 AND Y = 43 else "111111110000" when X = 61 AND Y = 43 else "111111110000" when X = 62 AND Y = 43 else "111111110000" when X = 63 AND Y = 43 else "111111110000" when X = 64 AND Y = 43 else "111111110000" when X = 65 AND Y = 43 else "111111110000" when X = 66 AND Y = 43 else "111111110000" when X = 67 AND Y = 43 else "111111110000" when X = 68 AND Y = 43 else "111111110000" when X = 0 AND Y = 44 else "111111110000" when X = 1 AND Y = 44 else "111111110000" when X = 2 AND Y = 44 else "111111110000" when X = 3 AND Y = 44 else "111111110000" when X = 4 AND Y = 44 else "111111110000" when X = 5 AND Y = 44 else "111111110000" when X = 6 AND Y = 44 else "111111110000" when X = 7 AND Y = 44 else "111111110000" when X = 8 AND Y = 44 else "111111110000" when X = 9 AND Y = 44 else "111111110000" when X = 10 AND Y = 44 else "111111110000" when X = 11 AND Y = 44 else "111111110000" when X = 12 AND Y = 44 else "111111110000" when X = 13 AND Y = 44 else "111111110000" when X = 14 AND Y = 44 else "111111110000" when X = 15 AND Y = 44 else "111111110000" when X = 16 AND Y = 44 else "111111110000" when X = 17 AND Y = 44 else "111111110000" when X = 18 AND Y = 44 else "111111110000" when X = 19 AND Y = 44 else "111111110000" when X = 20 AND Y = 44 else "111111110000" when X = 21 AND Y = 44 else "111111110000" when X = 22 AND Y = 44 else "111111110000" when X = 23 AND Y = 44 else "111111110000" when X = 24 AND Y = 44 else "111111110000" when X = 25 AND Y = 44 else "111111110000" when X = 26 AND Y = 44 else "111111110000" when X = 27 AND Y = 44 else "111111110000" when X = 28 AND Y = 44 else "111111110000" when X = 29 AND Y = 44 else "111111110000" when X = 30 AND Y = 44 else "111111110000" when X = 31 AND Y = 44 else "111111110000" when X = 32 AND Y = 44 else "111111110000" when X = 33 AND Y = 44 else "111111110000" when X = 34 AND Y = 44 else "111111110000" when X = 35 AND Y = 44 else "111111110000" when X = 36 AND Y = 44 else "111111110000" when X = 37 AND Y = 44 else "111111110000" when X = 38 AND Y = 44 else "111111110000" when X = 39 AND Y = 44 else "111111110000" when X = 40 AND Y = 44 else "111111110000" when X = 41 AND Y = 44 else "111111110000" when X = 42 AND Y = 44 else "111111110000" when X = 43 AND Y = 44 else "111111110000" when X = 44 AND Y = 44 else "111111110000" when X = 45 AND Y = 44 else "111111110000" when X = 46 AND Y = 44 else "111111110000" when X = 47 AND Y = 44 else "111111110000" when X = 48 AND Y = 44 else "111111110000" when X = 49 AND Y = 44 else "111111110000" when X = 50 AND Y = 44 else "111111110000" when X = 51 AND Y = 44 else "111111110000" when X = 52 AND Y = 44 else "111111110000" when X = 53 AND Y = 44 else "111111110000" when X = 54 AND Y = 44 else "111111110000" when X = 55 AND Y = 44 else "111111110000" when X = 56 AND Y = 44 else "111111110000" when X = 57 AND Y = 44 else "111111110000" when X = 58 AND Y = 44 else "111111110000" when X = 59 AND Y = 44 else "111111110000" when X = 60 AND Y = 44 else "111111110000" when X = 61 AND Y = 44 else "111111110000" when X = 62 AND Y = 44 else "111111110000" when X = 63 AND Y = 44 else "111111110000" when X = 64 AND Y = 44 else "111111110000" when X = 65 AND Y = 44 else "111111110000" when X = 66 AND Y = 44 else "111111110000" when X = 67 AND Y = 44 else "111111110000" when X = 68 AND Y = 44 else 
"000000000000"; -- should never get here
end rtl;
