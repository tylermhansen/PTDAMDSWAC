-- Tyler Hansen
-- CS232 Final Project
-- genSpriteROM.py
-- generates a ROM file in VHDL from a .ppm image

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity cloud is
port(
X	: in INTEGER RANGE 0 TO 1688;
Y	: in INTEGER RANGE 0 TO 1688;
data : out std_logic_vector (11 downto 0)
);

end entity;

architecture rtl of cloud is
begin
data <=
"000000000000" when X = 0 AND Y = 0 else
"000000000000" when X = 1 AND Y = 0 else
"000000000000" when X = 2 AND Y = 0 else
"000000000000" when X = 3 AND Y = 0 else
"000000000000" when X = 4 AND Y = 0 else
"000000000000" when X = 5 AND Y = 0 else
"000000000000" when X = 6 AND Y = 0 else
"000000000000" when X = 7 AND Y = 0 else
"000000000000" when X = 8 AND Y = 0 else
"000000000000" when X = 9 AND Y = 0 else
"000000000000" when X = 10 AND Y = 0 else
"000000000000" when X = 11 AND Y = 0 else
"000000000000" when X = 12 AND Y = 0 else
"000000000000" when X = 13 AND Y = 0 else
"000100010001" when X = 14 AND Y = 0 else
"001100110011" when X = 15 AND Y = 0 else
"001100110100" when X = 16 AND Y = 0 else
"010001000100" when X = 17 AND Y = 0 else
"110011001100" when X = 18 AND Y = 0 else
"111111111111" when X = 19 AND Y = 0 else
"111111111111" when X = 20 AND Y = 0 else
"111111111111" when X = 21 AND Y = 0 else
"111111111111" when X = 22 AND Y = 0 else
"111111111111" when X = 23 AND Y = 0 else
"111111111111" when X = 24 AND Y = 0 else
"111111111111" when X = 25 AND Y = 0 else
"111111111111" when X = 26 AND Y = 0 else
"111111111111" when X = 27 AND Y = 0 else
"111111111111" when X = 28 AND Y = 0 else
"111111111111" when X = 29 AND Y = 0 else
"111111111111" when X = 30 AND Y = 0 else
"111111111111" when X = 31 AND Y = 0 else
"101010101010" when X = 32 AND Y = 0 else
"001000100010" when X = 33 AND Y = 0 else
"000000000000" when X = 34 AND Y = 0 else
"000000000000" when X = 35 AND Y = 0 else
"000000000000" when X = 36 AND Y = 0 else
"000000000000" when X = 37 AND Y = 0 else
"000000000000" when X = 38 AND Y = 0 else
"000000000000" when X = 39 AND Y = 0 else
"000000000000" when X = 40 AND Y = 0 else
"000000000000" when X = 41 AND Y = 0 else
"000000000000" when X = 42 AND Y = 0 else
"000000000000" when X = 43 AND Y = 0 else
"000000000000" when X = 44 AND Y = 0 else
"000000000000" when X = 45 AND Y = 0 else
"000000000000" when X = 46 AND Y = 0 else
"000000000000" when X = 47 AND Y = 0 else
"000000000000" when X = 48 AND Y = 0 else
"000000000000" when X = 49 AND Y = 0 else
"000000000000" when X = 50 AND Y = 0 else
"000000000000" when X = 51 AND Y = 0 else
"000000000000" when X = 52 AND Y = 0 else
"000000000000" when X = 53 AND Y = 0 else
"000000000000" when X = 54 AND Y = 0 else
"000000000000" when X = 55 AND Y = 0 else
"000000000000" when X = 56 AND Y = 0 else
"000000000000" when X = 57 AND Y = 0 else
"000000000000" when X = 58 AND Y = 0 else
"000000000000" when X = 59 AND Y = 0 else
"000000000000" when X = 60 AND Y = 0 else
"000000000000" when X = 61 AND Y = 0 else
"000000000000" when X = 62 AND Y = 0 else
"000000000000" when X = 63 AND Y = 0 else
"000000000000" when X = 64 AND Y = 0 else
"000000000000" when X = 65 AND Y = 0 else
"000000000000" when X = 66 AND Y = 0 else
"000000000000" when X = 67 AND Y = 0 else
"000000000000" when X = 68 AND Y = 0 else
"000000000000" when X = 69 AND Y = 0 else
"000000000000" when X = 70 AND Y = 0 else
"000000000000" when X = 71 AND Y = 0 else
"000000000000" when X = 72 AND Y = 0 else
"000000000000" when X = 73 AND Y = 0 else
"000000000000" when X = 74 AND Y = 0 else
"000000000000" when X = 0 AND Y = 1 else
"000000000000" when X = 1 AND Y = 1 else
"000000000000" when X = 2 AND Y = 1 else
"000000000000" when X = 3 AND Y = 1 else
"000000000000" when X = 4 AND Y = 1 else
"000000000000" when X = 5 AND Y = 1 else
"000000000000" when X = 6 AND Y = 1 else
"000000000000" when X = 7 AND Y = 1 else
"000000000000" when X = 8 AND Y = 1 else
"000000000000" when X = 9 AND Y = 1 else
"000000000000" when X = 10 AND Y = 1 else
"000000000000" when X = 11 AND Y = 1 else
"000000000000" when X = 12 AND Y = 1 else
"000000000000" when X = 13 AND Y = 1 else
"010001000101" when X = 14 AND Y = 1 else
"101110111100" when X = 15 AND Y = 1 else
"110011001101" when X = 16 AND Y = 1 else
"110111011110" when X = 17 AND Y = 1 else
"111111111111" when X = 18 AND Y = 1 else
"111111111111" when X = 19 AND Y = 1 else
"111111111111" when X = 20 AND Y = 1 else
"111111111111" when X = 21 AND Y = 1 else
"111111111111" when X = 22 AND Y = 1 else
"111111111111" when X = 23 AND Y = 1 else
"111111111111" when X = 24 AND Y = 1 else
"111111111111" when X = 25 AND Y = 1 else
"111111111111" when X = 26 AND Y = 1 else
"111111111111" when X = 27 AND Y = 1 else
"111111111111" when X = 28 AND Y = 1 else
"111111111111" when X = 29 AND Y = 1 else
"111111111111" when X = 30 AND Y = 1 else
"111111111111" when X = 31 AND Y = 1 else
"111011101110" when X = 32 AND Y = 1 else
"101010101010" when X = 33 AND Y = 1 else
"000000000000" when X = 34 AND Y = 1 else
"000000000000" when X = 35 AND Y = 1 else
"000000000000" when X = 36 AND Y = 1 else
"000000000000" when X = 37 AND Y = 1 else
"000000000000" when X = 38 AND Y = 1 else
"000000000000" when X = 39 AND Y = 1 else
"000000000000" when X = 40 AND Y = 1 else
"000000000000" when X = 41 AND Y = 1 else
"000000000000" when X = 42 AND Y = 1 else
"000000000000" when X = 43 AND Y = 1 else
"000000000000" when X = 44 AND Y = 1 else
"000000000000" when X = 45 AND Y = 1 else
"000000000000" when X = 46 AND Y = 1 else
"000000000000" when X = 47 AND Y = 1 else
"000000000000" when X = 48 AND Y = 1 else
"000000000000" when X = 49 AND Y = 1 else
"000000000000" when X = 50 AND Y = 1 else
"000000000000" when X = 51 AND Y = 1 else
"000000000000" when X = 52 AND Y = 1 else
"000000000000" when X = 53 AND Y = 1 else
"000000000000" when X = 54 AND Y = 1 else
"000000000000" when X = 55 AND Y = 1 else
"000000000000" when X = 56 AND Y = 1 else
"000000000000" when X = 57 AND Y = 1 else
"000000000000" when X = 58 AND Y = 1 else
"000000000000" when X = 59 AND Y = 1 else
"000000000000" when X = 60 AND Y = 1 else
"000000000000" when X = 61 AND Y = 1 else
"000000000000" when X = 62 AND Y = 1 else
"000000000000" when X = 63 AND Y = 1 else
"000000000000" when X = 64 AND Y = 1 else
"000000000000" when X = 65 AND Y = 1 else
"000000000000" when X = 66 AND Y = 1 else
"000000000000" when X = 67 AND Y = 1 else
"000000000000" when X = 68 AND Y = 1 else
"000000000000" when X = 69 AND Y = 1 else
"000000000000" when X = 70 AND Y = 1 else
"000000000000" when X = 71 AND Y = 1 else
"000000000000" when X = 72 AND Y = 1 else
"000000000000" when X = 73 AND Y = 1 else
"000000000000" when X = 74 AND Y = 1 else
"000000000000" when X = 0 AND Y = 2 else
"000000000000" when X = 1 AND Y = 2 else
"000000000000" when X = 2 AND Y = 2 else
"000000000000" when X = 3 AND Y = 2 else
"000000000000" when X = 4 AND Y = 2 else
"000000000000" when X = 5 AND Y = 2 else
"000000000000" when X = 6 AND Y = 2 else
"000000000000" when X = 7 AND Y = 2 else
"000000000000" when X = 8 AND Y = 2 else
"000000000000" when X = 9 AND Y = 2 else
"000000000000" when X = 10 AND Y = 2 else
"000000000000" when X = 11 AND Y = 2 else
"000000000000" when X = 12 AND Y = 2 else
"010101010110" when X = 13 AND Y = 2 else
"101110111100" when X = 14 AND Y = 2 else
"110111011110" when X = 15 AND Y = 2 else
"111011101111" when X = 16 AND Y = 2 else
"111111111111" when X = 17 AND Y = 2 else
"111111111111" when X = 18 AND Y = 2 else
"111111111111" when X = 19 AND Y = 2 else
"111111111111" when X = 20 AND Y = 2 else
"111111111111" when X = 21 AND Y = 2 else
"111111111111" when X = 22 AND Y = 2 else
"111111111111" when X = 23 AND Y = 2 else
"111111111111" when X = 24 AND Y = 2 else
"111111111111" when X = 25 AND Y = 2 else
"111111111111" when X = 26 AND Y = 2 else
"111111111111" when X = 27 AND Y = 2 else
"111111111111" when X = 28 AND Y = 2 else
"111111111111" when X = 29 AND Y = 2 else
"111111111111" when X = 30 AND Y = 2 else
"111111111111" when X = 31 AND Y = 2 else
"111111111111" when X = 32 AND Y = 2 else
"111011101110" when X = 33 AND Y = 2 else
"101010101010" when X = 34 AND Y = 2 else
"000000000000" when X = 35 AND Y = 2 else
"000000000000" when X = 36 AND Y = 2 else
"000000000000" when X = 37 AND Y = 2 else
"000000000000" when X = 38 AND Y = 2 else
"000000000000" when X = 39 AND Y = 2 else
"000000000000" when X = 40 AND Y = 2 else
"000000000000" when X = 41 AND Y = 2 else
"000000000000" when X = 42 AND Y = 2 else
"000000000000" when X = 43 AND Y = 2 else
"000000000000" when X = 44 AND Y = 2 else
"000000000000" when X = 45 AND Y = 2 else
"000000000000" when X = 46 AND Y = 2 else
"000000000000" when X = 47 AND Y = 2 else
"000000000000" when X = 48 AND Y = 2 else
"000000000000" when X = 49 AND Y = 2 else
"000000000000" when X = 50 AND Y = 2 else
"000000000000" when X = 51 AND Y = 2 else
"000000000000" when X = 52 AND Y = 2 else
"000000000000" when X = 53 AND Y = 2 else
"000000000000" when X = 54 AND Y = 2 else
"000000000000" when X = 55 AND Y = 2 else
"000000000000" when X = 56 AND Y = 2 else
"000000000000" when X = 57 AND Y = 2 else
"000000000000" when X = 58 AND Y = 2 else
"000000000000" when X = 59 AND Y = 2 else
"000000000000" when X = 60 AND Y = 2 else
"000000000000" when X = 61 AND Y = 2 else
"000000000000" when X = 62 AND Y = 2 else
"000000000000" when X = 63 AND Y = 2 else
"000000000000" when X = 64 AND Y = 2 else
"000000000000" when X = 65 AND Y = 2 else
"000000000000" when X = 66 AND Y = 2 else
"000000000000" when X = 67 AND Y = 2 else
"000000000000" when X = 68 AND Y = 2 else
"000000000000" when X = 69 AND Y = 2 else
"000000000000" when X = 70 AND Y = 2 else
"000000000000" when X = 71 AND Y = 2 else
"000000000000" when X = 72 AND Y = 2 else
"000000000000" when X = 73 AND Y = 2 else
"000000000000" when X = 74 AND Y = 2 else
"000000000000" when X = 0 AND Y = 3 else
"000000000000" when X = 1 AND Y = 3 else
"000000000000" when X = 2 AND Y = 3 else
"000000000000" when X = 3 AND Y = 3 else
"000000000000" when X = 4 AND Y = 3 else
"000000000000" when X = 5 AND Y = 3 else
"000000000000" when X = 6 AND Y = 3 else
"000000000000" when X = 7 AND Y = 3 else
"000000000000" when X = 8 AND Y = 3 else
"000000000000" when X = 9 AND Y = 3 else
"000000000000" when X = 10 AND Y = 3 else
"011101111000" when X = 11 AND Y = 3 else
"101010101011" when X = 12 AND Y = 3 else
"101110111100" when X = 13 AND Y = 3 else
"110111011111" when X = 14 AND Y = 3 else
"111011101111" when X = 15 AND Y = 3 else
"111111111111" when X = 16 AND Y = 3 else
"111111111111" when X = 17 AND Y = 3 else
"111111111111" when X = 18 AND Y = 3 else
"111111111111" when X = 19 AND Y = 3 else
"111111111111" when X = 20 AND Y = 3 else
"111111111111" when X = 21 AND Y = 3 else
"111111111111" when X = 22 AND Y = 3 else
"111111111111" when X = 23 AND Y = 3 else
"111111111111" when X = 24 AND Y = 3 else
"111111111111" when X = 25 AND Y = 3 else
"111111111111" when X = 26 AND Y = 3 else
"111111111111" when X = 27 AND Y = 3 else
"111111111111" when X = 28 AND Y = 3 else
"111111111111" when X = 29 AND Y = 3 else
"111111111111" when X = 30 AND Y = 3 else
"111111111111" when X = 31 AND Y = 3 else
"111111111111" when X = 32 AND Y = 3 else
"111111111111" when X = 33 AND Y = 3 else
"111011101110" when X = 34 AND Y = 3 else
"101010101010" when X = 35 AND Y = 3 else
"001000100010" when X = 36 AND Y = 3 else
"000000000000" when X = 37 AND Y = 3 else
"000000000000" when X = 38 AND Y = 3 else
"000000000000" when X = 39 AND Y = 3 else
"000000000000" when X = 40 AND Y = 3 else
"000000000000" when X = 41 AND Y = 3 else
"000000000000" when X = 42 AND Y = 3 else
"000000000000" when X = 43 AND Y = 3 else
"000000000000" when X = 44 AND Y = 3 else
"000000000000" when X = 45 AND Y = 3 else
"000000000000" when X = 46 AND Y = 3 else
"000000000000" when X = 47 AND Y = 3 else
"000000000000" when X = 48 AND Y = 3 else
"000000000000" when X = 49 AND Y = 3 else
"000000000000" when X = 50 AND Y = 3 else
"000000000000" when X = 51 AND Y = 3 else
"000000000000" when X = 52 AND Y = 3 else
"000000000000" when X = 53 AND Y = 3 else
"000000000000" when X = 54 AND Y = 3 else
"000000000000" when X = 55 AND Y = 3 else
"000000000000" when X = 56 AND Y = 3 else
"000000000000" when X = 57 AND Y = 3 else
"000000000000" when X = 58 AND Y = 3 else
"000000000000" when X = 59 AND Y = 3 else
"000000000000" when X = 60 AND Y = 3 else
"000000000000" when X = 61 AND Y = 3 else
"000000000000" when X = 62 AND Y = 3 else
"000000000000" when X = 63 AND Y = 3 else
"000000000000" when X = 64 AND Y = 3 else
"000000000000" when X = 65 AND Y = 3 else
"000000000000" when X = 66 AND Y = 3 else
"000000000000" when X = 67 AND Y = 3 else
"000000000000" when X = 68 AND Y = 3 else
"000000000000" when X = 69 AND Y = 3 else
"000000000000" when X = 70 AND Y = 3 else
"000000000000" when X = 71 AND Y = 3 else
"000000000000" when X = 72 AND Y = 3 else
"000000000000" when X = 73 AND Y = 3 else
"000000000000" when X = 74 AND Y = 3 else
"000000000000" when X = 0 AND Y = 4 else
"000000000000" when X = 1 AND Y = 4 else
"000000000000" when X = 2 AND Y = 4 else
"000000000000" when X = 3 AND Y = 4 else
"000000000000" when X = 4 AND Y = 4 else
"000000000000" when X = 5 AND Y = 4 else
"000000000000" when X = 6 AND Y = 4 else
"000000000000" when X = 7 AND Y = 4 else
"000000000000" when X = 8 AND Y = 4 else
"000000000000" when X = 9 AND Y = 4 else
"010001000111" when X = 10 AND Y = 4 else
"100110101100" when X = 11 AND Y = 4 else
"110111011111" when X = 12 AND Y = 4 else
"110111011111" when X = 13 AND Y = 4 else
"111011101111" when X = 14 AND Y = 4 else
"111111111111" when X = 15 AND Y = 4 else
"111111111111" when X = 16 AND Y = 4 else
"111111111111" when X = 17 AND Y = 4 else
"111111111111" when X = 18 AND Y = 4 else
"111111111111" when X = 19 AND Y = 4 else
"111111111111" when X = 20 AND Y = 4 else
"111111111111" when X = 21 AND Y = 4 else
"111111111111" when X = 22 AND Y = 4 else
"111111111111" when X = 23 AND Y = 4 else
"111111111111" when X = 24 AND Y = 4 else
"111111111111" when X = 25 AND Y = 4 else
"111111111111" when X = 26 AND Y = 4 else
"111111111111" when X = 27 AND Y = 4 else
"111111111111" when X = 28 AND Y = 4 else
"111111111111" when X = 29 AND Y = 4 else
"111111111111" when X = 30 AND Y = 4 else
"111111111111" when X = 31 AND Y = 4 else
"111111111111" when X = 32 AND Y = 4 else
"111111111111" when X = 33 AND Y = 4 else
"111111111111" when X = 34 AND Y = 4 else
"110111011101" when X = 35 AND Y = 4 else
"000100010001" when X = 36 AND Y = 4 else
"000000000000" when X = 37 AND Y = 4 else
"000000000000" when X = 38 AND Y = 4 else
"000000000000" when X = 39 AND Y = 4 else
"000000000000" when X = 40 AND Y = 4 else
"000000000000" when X = 41 AND Y = 4 else
"000000000000" when X = 42 AND Y = 4 else
"000000000000" when X = 43 AND Y = 4 else
"000000000000" when X = 44 AND Y = 4 else
"000000000000" when X = 45 AND Y = 4 else
"000000000000" when X = 46 AND Y = 4 else
"000000000000" when X = 47 AND Y = 4 else
"000000000000" when X = 48 AND Y = 4 else
"000000000000" when X = 49 AND Y = 4 else
"000000000000" when X = 50 AND Y = 4 else
"000000000000" when X = 51 AND Y = 4 else
"000000000000" when X = 52 AND Y = 4 else
"000000000000" when X = 53 AND Y = 4 else
"000000000000" when X = 54 AND Y = 4 else
"000000000000" when X = 55 AND Y = 4 else
"000000000000" when X = 56 AND Y = 4 else
"000000000000" when X = 57 AND Y = 4 else
"000000000000" when X = 58 AND Y = 4 else
"000000000000" when X = 59 AND Y = 4 else
"000000000000" when X = 60 AND Y = 4 else
"000000000000" when X = 61 AND Y = 4 else
"000000000000" when X = 62 AND Y = 4 else
"000000000000" when X = 63 AND Y = 4 else
"000000000000" when X = 64 AND Y = 4 else
"000000000000" when X = 65 AND Y = 4 else
"000000000000" when X = 66 AND Y = 4 else
"000000000000" when X = 67 AND Y = 4 else
"000000000000" when X = 68 AND Y = 4 else
"000000000000" when X = 69 AND Y = 4 else
"000000000000" when X = 70 AND Y = 4 else
"000000000000" when X = 71 AND Y = 4 else
"000000000000" when X = 72 AND Y = 4 else
"000000000000" when X = 73 AND Y = 4 else
"000000000000" when X = 74 AND Y = 4 else
"000000000000" when X = 0 AND Y = 5 else
"000000000000" when X = 1 AND Y = 5 else
"000000000000" when X = 2 AND Y = 5 else
"000000000000" when X = 3 AND Y = 5 else
"000000000000" when X = 4 AND Y = 5 else
"000000000000" when X = 5 AND Y = 5 else
"000000000000" when X = 6 AND Y = 5 else
"000000000000" when X = 7 AND Y = 5 else
"000000000000" when X = 8 AND Y = 5 else
"000000000000" when X = 9 AND Y = 5 else
"011001111010" when X = 10 AND Y = 5 else
"101010111110" when X = 11 AND Y = 5 else
"110111011111" when X = 12 AND Y = 5 else
"110111101111" when X = 13 AND Y = 5 else
"111111111111" when X = 14 AND Y = 5 else
"111111111111" when X = 15 AND Y = 5 else
"111111111111" when X = 16 AND Y = 5 else
"111111111111" when X = 17 AND Y = 5 else
"111111111111" when X = 18 AND Y = 5 else
"111111111111" when X = 19 AND Y = 5 else
"111111111111" when X = 20 AND Y = 5 else
"111111111111" when X = 21 AND Y = 5 else
"111111111111" when X = 22 AND Y = 5 else
"111111111111" when X = 23 AND Y = 5 else
"111111111111" when X = 24 AND Y = 5 else
"111111111111" when X = 25 AND Y = 5 else
"111111111111" when X = 26 AND Y = 5 else
"111111111111" when X = 27 AND Y = 5 else
"111111111111" when X = 28 AND Y = 5 else
"111111111111" when X = 29 AND Y = 5 else
"111111111111" when X = 30 AND Y = 5 else
"111111111111" when X = 31 AND Y = 5 else
"111111111111" when X = 32 AND Y = 5 else
"111111111111" when X = 33 AND Y = 5 else
"111111111111" when X = 34 AND Y = 5 else
"111011101110" when X = 35 AND Y = 5 else
"100010001000" when X = 36 AND Y = 5 else
"000100010001" when X = 37 AND Y = 5 else
"000000000000" when X = 38 AND Y = 5 else
"000000000000" when X = 39 AND Y = 5 else
"000000000000" when X = 40 AND Y = 5 else
"000000000000" when X = 41 AND Y = 5 else
"000000000000" when X = 42 AND Y = 5 else
"000000000000" when X = 43 AND Y = 5 else
"000000000000" when X = 44 AND Y = 5 else
"000000000000" when X = 45 AND Y = 5 else
"000000000000" when X = 46 AND Y = 5 else
"000000000000" when X = 47 AND Y = 5 else
"000000000000" when X = 48 AND Y = 5 else
"000000000000" when X = 49 AND Y = 5 else
"000000000000" when X = 50 AND Y = 5 else
"000000000000" when X = 51 AND Y = 5 else
"000000000000" when X = 52 AND Y = 5 else
"000000000000" when X = 53 AND Y = 5 else
"011101110111" when X = 54 AND Y = 5 else
"100110011001" when X = 55 AND Y = 5 else
"100110011001" when X = 56 AND Y = 5 else
"100010001001" when X = 57 AND Y = 5 else
"011101111000" when X = 58 AND Y = 5 else
"011101111000" when X = 59 AND Y = 5 else
"011101111000" when X = 60 AND Y = 5 else
"011101111000" when X = 61 AND Y = 5 else
"010001000101" when X = 62 AND Y = 5 else
"000000000000" when X = 63 AND Y = 5 else
"000000000000" when X = 64 AND Y = 5 else
"000000000000" when X = 65 AND Y = 5 else
"000000000000" when X = 66 AND Y = 5 else
"000000000000" when X = 67 AND Y = 5 else
"000000000000" when X = 68 AND Y = 5 else
"000000000000" when X = 69 AND Y = 5 else
"000000000000" when X = 70 AND Y = 5 else
"000000000000" when X = 71 AND Y = 5 else
"000000000000" when X = 72 AND Y = 5 else
"000000000000" when X = 73 AND Y = 5 else
"000000000000" when X = 74 AND Y = 5 else
"000000000000" when X = 0 AND Y = 6 else
"000000000000" when X = 1 AND Y = 6 else
"000000000000" when X = 2 AND Y = 6 else
"000000000000" when X = 3 AND Y = 6 else
"000000000000" when X = 4 AND Y = 6 else
"000000000000" when X = 5 AND Y = 6 else
"000000000000" when X = 6 AND Y = 6 else
"000000000000" when X = 7 AND Y = 6 else
"000000000000" when X = 8 AND Y = 6 else
"000000000000" when X = 9 AND Y = 6 else
"011001111010" when X = 10 AND Y = 6 else
"101010111110" when X = 11 AND Y = 6 else
"110111011111" when X = 12 AND Y = 6 else
"110111101111" when X = 13 AND Y = 6 else
"111111111111" when X = 14 AND Y = 6 else
"111111111111" when X = 15 AND Y = 6 else
"111111111111" when X = 16 AND Y = 6 else
"111111111111" when X = 17 AND Y = 6 else
"111111111111" when X = 18 AND Y = 6 else
"111111111111" when X = 19 AND Y = 6 else
"111111111111" when X = 20 AND Y = 6 else
"111111111111" when X = 21 AND Y = 6 else
"111111111111" when X = 22 AND Y = 6 else
"111111111111" when X = 23 AND Y = 6 else
"111111111111" when X = 24 AND Y = 6 else
"111111111111" when X = 25 AND Y = 6 else
"111111111111" when X = 26 AND Y = 6 else
"111111111111" when X = 27 AND Y = 6 else
"111111111111" when X = 28 AND Y = 6 else
"111111111111" when X = 29 AND Y = 6 else
"111111111111" when X = 30 AND Y = 6 else
"111111111111" when X = 31 AND Y = 6 else
"111111111111" when X = 32 AND Y = 6 else
"111111111111" when X = 33 AND Y = 6 else
"111111111111" when X = 34 AND Y = 6 else
"111111111111" when X = 35 AND Y = 6 else
"111011101110" when X = 36 AND Y = 6 else
"100010001000" when X = 37 AND Y = 6 else
"011101110111" when X = 38 AND Y = 6 else
"011101110111" when X = 39 AND Y = 6 else
"011101110111" when X = 40 AND Y = 6 else
"011101110111" when X = 41 AND Y = 6 else
"011101110111" when X = 42 AND Y = 6 else
"011001100110" when X = 43 AND Y = 6 else
"000000000000" when X = 44 AND Y = 6 else
"000000000000" when X = 45 AND Y = 6 else
"000000000000" when X = 46 AND Y = 6 else
"000000000000" when X = 47 AND Y = 6 else
"000000000000" when X = 48 AND Y = 6 else
"000000000000" when X = 49 AND Y = 6 else
"000000000000" when X = 50 AND Y = 6 else
"001000100010" when X = 51 AND Y = 6 else
"011101110111" when X = 52 AND Y = 6 else
"011101110111" when X = 53 AND Y = 6 else
"111011101110" when X = 54 AND Y = 6 else
"111111111111" when X = 55 AND Y = 6 else
"111111111111" when X = 56 AND Y = 6 else
"111111111111" when X = 57 AND Y = 6 else
"110111011111" when X = 58 AND Y = 6 else
"110111011110" when X = 59 AND Y = 6 else
"110111011110" when X = 60 AND Y = 6 else
"110111011110" when X = 61 AND Y = 6 else
"100110011010" when X = 62 AND Y = 6 else
"010001000100" when X = 63 AND Y = 6 else
"000000000000" when X = 64 AND Y = 6 else
"000000000000" when X = 65 AND Y = 6 else
"000000000000" when X = 66 AND Y = 6 else
"000000000000" when X = 67 AND Y = 6 else
"000000000000" when X = 68 AND Y = 6 else
"000000000000" when X = 69 AND Y = 6 else
"000000000000" when X = 70 AND Y = 6 else
"000000000000" when X = 71 AND Y = 6 else
"000000000000" when X = 72 AND Y = 6 else
"000000000000" when X = 73 AND Y = 6 else
"000000000000" when X = 74 AND Y = 6 else
"000000000000" when X = 0 AND Y = 7 else
"000000000000" when X = 1 AND Y = 7 else
"000000000000" when X = 2 AND Y = 7 else
"000000000000" when X = 3 AND Y = 7 else
"000000000000" when X = 4 AND Y = 7 else
"000000000000" when X = 5 AND Y = 7 else
"000000000000" when X = 6 AND Y = 7 else
"000000000000" when X = 7 AND Y = 7 else
"000000000000" when X = 8 AND Y = 7 else
"000000000000" when X = 9 AND Y = 7 else
"011001111010" when X = 10 AND Y = 7 else
"101010111110" when X = 11 AND Y = 7 else
"110111011111" when X = 12 AND Y = 7 else
"110111101111" when X = 13 AND Y = 7 else
"111111111111" when X = 14 AND Y = 7 else
"111111111111" when X = 15 AND Y = 7 else
"111111111111" when X = 16 AND Y = 7 else
"111111111111" when X = 17 AND Y = 7 else
"111111111111" when X = 18 AND Y = 7 else
"111111111111" when X = 19 AND Y = 7 else
"111111111111" when X = 20 AND Y = 7 else
"111111111111" when X = 21 AND Y = 7 else
"111111111111" when X = 22 AND Y = 7 else
"111111111111" when X = 23 AND Y = 7 else
"111111111111" when X = 24 AND Y = 7 else
"111111111111" when X = 25 AND Y = 7 else
"111111111111" when X = 26 AND Y = 7 else
"111111111111" when X = 27 AND Y = 7 else
"111111111111" when X = 28 AND Y = 7 else
"111111111111" when X = 29 AND Y = 7 else
"111111111111" when X = 30 AND Y = 7 else
"111111111111" when X = 31 AND Y = 7 else
"111111111111" when X = 32 AND Y = 7 else
"111111111111" when X = 33 AND Y = 7 else
"111111111111" when X = 34 AND Y = 7 else
"111111111111" when X = 35 AND Y = 7 else
"111111111111" when X = 36 AND Y = 7 else
"111111111111" when X = 37 AND Y = 7 else
"111111111111" when X = 38 AND Y = 7 else
"111111111111" when X = 39 AND Y = 7 else
"111111111111" when X = 40 AND Y = 7 else
"111111111111" when X = 41 AND Y = 7 else
"111111111111" when X = 42 AND Y = 7 else
"111011101110" when X = 43 AND Y = 7 else
"011001100110" when X = 44 AND Y = 7 else
"010101010101" when X = 45 AND Y = 7 else
"001000100010" when X = 46 AND Y = 7 else
"000000000000" when X = 47 AND Y = 7 else
"000000000000" when X = 48 AND Y = 7 else
"001100110011" when X = 49 AND Y = 7 else
"010101010101" when X = 50 AND Y = 7 else
"100010001000" when X = 51 AND Y = 7 else
"111011101110" when X = 52 AND Y = 7 else
"111111111111" when X = 53 AND Y = 7 else
"111111111111" when X = 54 AND Y = 7 else
"111111111111" when X = 55 AND Y = 7 else
"111111111111" when X = 56 AND Y = 7 else
"111111111111" when X = 57 AND Y = 7 else
"111111111111" when X = 58 AND Y = 7 else
"110111101111" when X = 59 AND Y = 7 else
"110111011111" when X = 60 AND Y = 7 else
"110111011111" when X = 61 AND Y = 7 else
"110111011110" when X = 62 AND Y = 7 else
"100110011010" when X = 63 AND Y = 7 else
"001100110100" when X = 64 AND Y = 7 else
"000000000000" when X = 65 AND Y = 7 else
"000000000000" when X = 66 AND Y = 7 else
"000000000000" when X = 67 AND Y = 7 else
"000000000000" when X = 68 AND Y = 7 else
"000000000000" when X = 69 AND Y = 7 else
"000000000000" when X = 70 AND Y = 7 else
"000000000000" when X = 71 AND Y = 7 else
"000000000000" when X = 72 AND Y = 7 else
"000000000000" when X = 73 AND Y = 7 else
"000000000000" when X = 74 AND Y = 7 else
"000000000000" when X = 0 AND Y = 8 else
"000000000000" when X = 1 AND Y = 8 else
"000000000000" when X = 2 AND Y = 8 else
"000000000000" when X = 3 AND Y = 8 else
"000000000000" when X = 4 AND Y = 8 else
"000000000000" when X = 5 AND Y = 8 else
"000000000000" when X = 6 AND Y = 8 else
"000000000000" when X = 7 AND Y = 8 else
"000000000000" when X = 8 AND Y = 8 else
"000000000000" when X = 9 AND Y = 8 else
"011001111010" when X = 10 AND Y = 8 else
"101010111110" when X = 11 AND Y = 8 else
"110111011111" when X = 12 AND Y = 8 else
"110111101111" when X = 13 AND Y = 8 else
"111111111111" when X = 14 AND Y = 8 else
"111111111111" when X = 15 AND Y = 8 else
"111111111111" when X = 16 AND Y = 8 else
"111111111111" when X = 17 AND Y = 8 else
"111111111111" when X = 18 AND Y = 8 else
"111111111111" when X = 19 AND Y = 8 else
"111111111111" when X = 20 AND Y = 8 else
"111111111111" when X = 21 AND Y = 8 else
"111111111111" when X = 22 AND Y = 8 else
"111111111111" when X = 23 AND Y = 8 else
"111111111111" when X = 24 AND Y = 8 else
"111111111111" when X = 25 AND Y = 8 else
"111111111111" when X = 26 AND Y = 8 else
"111111111111" when X = 27 AND Y = 8 else
"111111111111" when X = 28 AND Y = 8 else
"111111111111" when X = 29 AND Y = 8 else
"111111111111" when X = 30 AND Y = 8 else
"111111111111" when X = 31 AND Y = 8 else
"111111111111" when X = 32 AND Y = 8 else
"111111111111" when X = 33 AND Y = 8 else
"111111111111" when X = 34 AND Y = 8 else
"111111111111" when X = 35 AND Y = 8 else
"111111111111" when X = 36 AND Y = 8 else
"111111111111" when X = 37 AND Y = 8 else
"111111111111" when X = 38 AND Y = 8 else
"111111111111" when X = 39 AND Y = 8 else
"111111111111" when X = 40 AND Y = 8 else
"111111111111" when X = 41 AND Y = 8 else
"111111111111" when X = 42 AND Y = 8 else
"111111111111" when X = 43 AND Y = 8 else
"111011101110" when X = 44 AND Y = 8 else
"111011101110" when X = 45 AND Y = 8 else
"100010001000" when X = 46 AND Y = 8 else
"001100110011" when X = 47 AND Y = 8 else
"001100110011" when X = 48 AND Y = 8 else
"101010101010" when X = 49 AND Y = 8 else
"111011101110" when X = 50 AND Y = 8 else
"111111111111" when X = 51 AND Y = 8 else
"111111111111" when X = 52 AND Y = 8 else
"111111111111" when X = 53 AND Y = 8 else
"111111111111" when X = 54 AND Y = 8 else
"111111111111" when X = 55 AND Y = 8 else
"111111111111" when X = 56 AND Y = 8 else
"111111111111" when X = 57 AND Y = 8 else
"111111111111" when X = 58 AND Y = 8 else
"111111111111" when X = 59 AND Y = 8 else
"110111101111" when X = 60 AND Y = 8 else
"110111011111" when X = 61 AND Y = 8 else
"110111011111" when X = 62 AND Y = 8 else
"110011011110" when X = 63 AND Y = 8 else
"100110101011" when X = 64 AND Y = 8 else
"000000000000" when X = 65 AND Y = 8 else
"000000000000" when X = 66 AND Y = 8 else
"000000000000" when X = 67 AND Y = 8 else
"000000000000" when X = 68 AND Y = 8 else
"000000000000" when X = 69 AND Y = 8 else
"000000000000" when X = 70 AND Y = 8 else
"000000000000" when X = 71 AND Y = 8 else
"000000000000" when X = 72 AND Y = 8 else
"000000000000" when X = 73 AND Y = 8 else
"000000000000" when X = 74 AND Y = 8 else
"000000000000" when X = 0 AND Y = 9 else
"000000000000" when X = 1 AND Y = 9 else
"000000000000" when X = 2 AND Y = 9 else
"000000000000" when X = 3 AND Y = 9 else
"000000000000" when X = 4 AND Y = 9 else
"000000000000" when X = 5 AND Y = 9 else
"000000000000" when X = 6 AND Y = 9 else
"000000000000" when X = 7 AND Y = 9 else
"000000000000" when X = 8 AND Y = 9 else
"000000000000" when X = 9 AND Y = 9 else
"011001111010" when X = 10 AND Y = 9 else
"101010111110" when X = 11 AND Y = 9 else
"110111011111" when X = 12 AND Y = 9 else
"110111101111" when X = 13 AND Y = 9 else
"111111111111" when X = 14 AND Y = 9 else
"111111111111" when X = 15 AND Y = 9 else
"111111111111" when X = 16 AND Y = 9 else
"111111111111" when X = 17 AND Y = 9 else
"111111111111" when X = 18 AND Y = 9 else
"111111111111" when X = 19 AND Y = 9 else
"111111111111" when X = 20 AND Y = 9 else
"111111111111" when X = 21 AND Y = 9 else
"111111111111" when X = 22 AND Y = 9 else
"111111111111" when X = 23 AND Y = 9 else
"111111111111" when X = 24 AND Y = 9 else
"111111111111" when X = 25 AND Y = 9 else
"111111111111" when X = 26 AND Y = 9 else
"111111111111" when X = 27 AND Y = 9 else
"111111111111" when X = 28 AND Y = 9 else
"111111111111" when X = 29 AND Y = 9 else
"111111111111" when X = 30 AND Y = 9 else
"111111111111" when X = 31 AND Y = 9 else
"111111111111" when X = 32 AND Y = 9 else
"111111111111" when X = 33 AND Y = 9 else
"111111111111" when X = 34 AND Y = 9 else
"111111111111" when X = 35 AND Y = 9 else
"111111111111" when X = 36 AND Y = 9 else
"111111111111" when X = 37 AND Y = 9 else
"111111111111" when X = 38 AND Y = 9 else
"111111111111" when X = 39 AND Y = 9 else
"111111111111" when X = 40 AND Y = 9 else
"111111111111" when X = 41 AND Y = 9 else
"111111111111" when X = 42 AND Y = 9 else
"111111111111" when X = 43 AND Y = 9 else
"111111111111" when X = 44 AND Y = 9 else
"111111111111" when X = 45 AND Y = 9 else
"111011101110" when X = 46 AND Y = 9 else
"111011101110" when X = 47 AND Y = 9 else
"111011101110" when X = 48 AND Y = 9 else
"111011101110" when X = 49 AND Y = 9 else
"111111111111" when X = 50 AND Y = 9 else
"111111111111" when X = 51 AND Y = 9 else
"111111111111" when X = 52 AND Y = 9 else
"111111111111" when X = 53 AND Y = 9 else
"111111111111" when X = 54 AND Y = 9 else
"111111111111" when X = 55 AND Y = 9 else
"111111111111" when X = 56 AND Y = 9 else
"111111111111" when X = 57 AND Y = 9 else
"111111111111" when X = 58 AND Y = 9 else
"111111111111" when X = 59 AND Y = 9 else
"111111111111" when X = 60 AND Y = 9 else
"110111101111" when X = 61 AND Y = 9 else
"110111011111" when X = 62 AND Y = 9 else
"110111011111" when X = 63 AND Y = 9 else
"101010101100" when X = 64 AND Y = 9 else
"000000000000" when X = 65 AND Y = 9 else
"000000000000" when X = 66 AND Y = 9 else
"000000000000" when X = 67 AND Y = 9 else
"000000000000" when X = 68 AND Y = 9 else
"000000000000" when X = 69 AND Y = 9 else
"000000000000" when X = 70 AND Y = 9 else
"000000000000" when X = 71 AND Y = 9 else
"000000000000" when X = 72 AND Y = 9 else
"000000000000" when X = 73 AND Y = 9 else
"000000000000" when X = 74 AND Y = 9 else
"000000000000" when X = 0 AND Y = 10 else
"000000000000" when X = 1 AND Y = 10 else
"000000000000" when X = 2 AND Y = 10 else
"000000000000" when X = 3 AND Y = 10 else
"000000000000" when X = 4 AND Y = 10 else
"000000000000" when X = 5 AND Y = 10 else
"000000000000" when X = 6 AND Y = 10 else
"000000000000" when X = 7 AND Y = 10 else
"000000000000" when X = 8 AND Y = 10 else
"000000000000" when X = 9 AND Y = 10 else
"011001111010" when X = 10 AND Y = 10 else
"101010111110" when X = 11 AND Y = 10 else
"110111011111" when X = 12 AND Y = 10 else
"110111101111" when X = 13 AND Y = 10 else
"111111111111" when X = 14 AND Y = 10 else
"111111111111" when X = 15 AND Y = 10 else
"111111111111" when X = 16 AND Y = 10 else
"111111111111" when X = 17 AND Y = 10 else
"111111111111" when X = 18 AND Y = 10 else
"111111111111" when X = 19 AND Y = 10 else
"111111111111" when X = 20 AND Y = 10 else
"111111111111" when X = 21 AND Y = 10 else
"111111111111" when X = 22 AND Y = 10 else
"111111111111" when X = 23 AND Y = 10 else
"111111111111" when X = 24 AND Y = 10 else
"111111111111" when X = 25 AND Y = 10 else
"111111111111" when X = 26 AND Y = 10 else
"111111111111" when X = 27 AND Y = 10 else
"111111111111" when X = 28 AND Y = 10 else
"111111111111" when X = 29 AND Y = 10 else
"111111111111" when X = 30 AND Y = 10 else
"111111111111" when X = 31 AND Y = 10 else
"111111111111" when X = 32 AND Y = 10 else
"111111111111" when X = 33 AND Y = 10 else
"111111111111" when X = 34 AND Y = 10 else
"111111111111" when X = 35 AND Y = 10 else
"111111111111" when X = 36 AND Y = 10 else
"111111111111" when X = 37 AND Y = 10 else
"111111111111" when X = 38 AND Y = 10 else
"111111111111" when X = 39 AND Y = 10 else
"111111111111" when X = 40 AND Y = 10 else
"111111111111" when X = 41 AND Y = 10 else
"111111111111" when X = 42 AND Y = 10 else
"111111111111" when X = 43 AND Y = 10 else
"111111111111" when X = 44 AND Y = 10 else
"111111111111" when X = 45 AND Y = 10 else
"111111111111" when X = 46 AND Y = 10 else
"111111111111" when X = 47 AND Y = 10 else
"111111111111" when X = 48 AND Y = 10 else
"111111111111" when X = 49 AND Y = 10 else
"111111111111" when X = 50 AND Y = 10 else
"111111111111" when X = 51 AND Y = 10 else
"111111111111" when X = 52 AND Y = 10 else
"111111111111" when X = 53 AND Y = 10 else
"111111111111" when X = 54 AND Y = 10 else
"111111111111" when X = 55 AND Y = 10 else
"111111111111" when X = 56 AND Y = 10 else
"111111111111" when X = 57 AND Y = 10 else
"111111111111" when X = 58 AND Y = 10 else
"111111111111" when X = 59 AND Y = 10 else
"111111111111" when X = 60 AND Y = 10 else
"110111101111" when X = 61 AND Y = 10 else
"110111011111" when X = 62 AND Y = 10 else
"110111011111" when X = 63 AND Y = 10 else
"101010101100" when X = 64 AND Y = 10 else
"000000000000" when X = 65 AND Y = 10 else
"000000000000" when X = 66 AND Y = 10 else
"000000000000" when X = 67 AND Y = 10 else
"000000000000" when X = 68 AND Y = 10 else
"000000000000" when X = 69 AND Y = 10 else
"000000000000" when X = 70 AND Y = 10 else
"000000000000" when X = 71 AND Y = 10 else
"000000000000" when X = 72 AND Y = 10 else
"000000000000" when X = 73 AND Y = 10 else
"000000000000" when X = 74 AND Y = 10 else
"000000000000" when X = 0 AND Y = 11 else
"000000000000" when X = 1 AND Y = 11 else
"000000000000" when X = 2 AND Y = 11 else
"000000000000" when X = 3 AND Y = 11 else
"000000000000" when X = 4 AND Y = 11 else
"000000000000" when X = 5 AND Y = 11 else
"000000000000" when X = 6 AND Y = 11 else
"000100010010" when X = 7 AND Y = 11 else
"010101101001" when X = 8 AND Y = 11 else
"010101101010" when X = 9 AND Y = 11 else
"100110011100" when X = 10 AND Y = 11 else
"110011001110" when X = 11 AND Y = 11 else
"110111011111" when X = 12 AND Y = 11 else
"110111011111" when X = 13 AND Y = 11 else
"111011101111" when X = 14 AND Y = 11 else
"111011101111" when X = 15 AND Y = 11 else
"111111111111" when X = 16 AND Y = 11 else
"111111111111" when X = 17 AND Y = 11 else
"111111111111" when X = 18 AND Y = 11 else
"111111111111" when X = 19 AND Y = 11 else
"111111111111" when X = 20 AND Y = 11 else
"111111111111" when X = 21 AND Y = 11 else
"111111111111" when X = 22 AND Y = 11 else
"111111111111" when X = 23 AND Y = 11 else
"111111111111" when X = 24 AND Y = 11 else
"111111111111" when X = 25 AND Y = 11 else
"111111111111" when X = 26 AND Y = 11 else
"111111111111" when X = 27 AND Y = 11 else
"111111111111" when X = 28 AND Y = 11 else
"111111111111" when X = 29 AND Y = 11 else
"111111111111" when X = 30 AND Y = 11 else
"111111111111" when X = 31 AND Y = 11 else
"111111111111" when X = 32 AND Y = 11 else
"111111111111" when X = 33 AND Y = 11 else
"111111111111" when X = 34 AND Y = 11 else
"111111111111" when X = 35 AND Y = 11 else
"111111111111" when X = 36 AND Y = 11 else
"111111111111" when X = 37 AND Y = 11 else
"111111111111" when X = 38 AND Y = 11 else
"111111111111" when X = 39 AND Y = 11 else
"111111111111" when X = 40 AND Y = 11 else
"111111111111" when X = 41 AND Y = 11 else
"111111111111" when X = 42 AND Y = 11 else
"111111111111" when X = 43 AND Y = 11 else
"111111111111" when X = 44 AND Y = 11 else
"111111111111" when X = 45 AND Y = 11 else
"111111111111" when X = 46 AND Y = 11 else
"111111111111" when X = 47 AND Y = 11 else
"111111111111" when X = 48 AND Y = 11 else
"111111111111" when X = 49 AND Y = 11 else
"111111111111" when X = 50 AND Y = 11 else
"111111111111" when X = 51 AND Y = 11 else
"111111111111" when X = 52 AND Y = 11 else
"111111111111" when X = 53 AND Y = 11 else
"111111111111" when X = 54 AND Y = 11 else
"111111111111" when X = 55 AND Y = 11 else
"111111111111" when X = 56 AND Y = 11 else
"111111111111" when X = 57 AND Y = 11 else
"111111111111" when X = 58 AND Y = 11 else
"111111111111" when X = 59 AND Y = 11 else
"111111111111" when X = 60 AND Y = 11 else
"110111101111" when X = 61 AND Y = 11 else
"110111011111" when X = 62 AND Y = 11 else
"110111011111" when X = 63 AND Y = 11 else
"101010101100" when X = 64 AND Y = 11 else
"000000000000" when X = 65 AND Y = 11 else
"000000000000" when X = 66 AND Y = 11 else
"000000000000" when X = 67 AND Y = 11 else
"000000000000" when X = 68 AND Y = 11 else
"000000000000" when X = 69 AND Y = 11 else
"000000000000" when X = 70 AND Y = 11 else
"000000000000" when X = 71 AND Y = 11 else
"000000000000" when X = 72 AND Y = 11 else
"000000000000" when X = 73 AND Y = 11 else
"000000000000" when X = 74 AND Y = 11 else
"000000000000" when X = 0 AND Y = 12 else
"000000000000" when X = 1 AND Y = 12 else
"000000000000" when X = 2 AND Y = 12 else
"000000000000" when X = 3 AND Y = 12 else
"000000000000" when X = 4 AND Y = 12 else
"000000000000" when X = 5 AND Y = 12 else
"000100100011" when X = 6 AND Y = 12 else
"010101101001" when X = 7 AND Y = 12 else
"011110001101" when X = 8 AND Y = 12 else
"100110101110" when X = 9 AND Y = 12 else
"110011001110" when X = 10 AND Y = 12 else
"110111011111" when X = 11 AND Y = 12 else
"110111011111" when X = 12 AND Y = 12 else
"110111011111" when X = 13 AND Y = 12 else
"110111011111" when X = 14 AND Y = 12 else
"110111011111" when X = 15 AND Y = 12 else
"111011101111" when X = 16 AND Y = 12 else
"111011111111" when X = 17 AND Y = 12 else
"111011111111" when X = 18 AND Y = 12 else
"111011111111" when X = 19 AND Y = 12 else
"111011111111" when X = 20 AND Y = 12 else
"111111111111" when X = 21 AND Y = 12 else
"111111111111" when X = 22 AND Y = 12 else
"111111111111" when X = 23 AND Y = 12 else
"111111111111" when X = 24 AND Y = 12 else
"111111111111" when X = 25 AND Y = 12 else
"111111111111" when X = 26 AND Y = 12 else
"111111111111" when X = 27 AND Y = 12 else
"111111111111" when X = 28 AND Y = 12 else
"111111111111" when X = 29 AND Y = 12 else
"111111111111" when X = 30 AND Y = 12 else
"111111111111" when X = 31 AND Y = 12 else
"111111111111" when X = 32 AND Y = 12 else
"111111111111" when X = 33 AND Y = 12 else
"111111111111" when X = 34 AND Y = 12 else
"111111111111" when X = 35 AND Y = 12 else
"111111111111" when X = 36 AND Y = 12 else
"111111111111" when X = 37 AND Y = 12 else
"111111111111" when X = 38 AND Y = 12 else
"111111111111" when X = 39 AND Y = 12 else
"111111111111" when X = 40 AND Y = 12 else
"111111111111" when X = 41 AND Y = 12 else
"111111111111" when X = 42 AND Y = 12 else
"111111111111" when X = 43 AND Y = 12 else
"111111111111" when X = 44 AND Y = 12 else
"111111111111" when X = 45 AND Y = 12 else
"111111111111" when X = 46 AND Y = 12 else
"111111111111" when X = 47 AND Y = 12 else
"111111111111" when X = 48 AND Y = 12 else
"111111111111" when X = 49 AND Y = 12 else
"111111111111" when X = 50 AND Y = 12 else
"111111111111" when X = 51 AND Y = 12 else
"111111111111" when X = 52 AND Y = 12 else
"111111111111" when X = 53 AND Y = 12 else
"111111111111" when X = 54 AND Y = 12 else
"111111111111" when X = 55 AND Y = 12 else
"111111111111" when X = 56 AND Y = 12 else
"111111111111" when X = 57 AND Y = 12 else
"111111111111" when X = 58 AND Y = 12 else
"111111111111" when X = 59 AND Y = 12 else
"111111111111" when X = 60 AND Y = 12 else
"110111101111" when X = 61 AND Y = 12 else
"110111011111" when X = 62 AND Y = 12 else
"110111011111" when X = 63 AND Y = 12 else
"101010101100" when X = 64 AND Y = 12 else
"000000000000" when X = 65 AND Y = 12 else
"000000000000" when X = 66 AND Y = 12 else
"000000000000" when X = 67 AND Y = 12 else
"000000000000" when X = 68 AND Y = 12 else
"000000000000" when X = 69 AND Y = 12 else
"000000000000" when X = 70 AND Y = 12 else
"000000000000" when X = 71 AND Y = 12 else
"000000000000" when X = 72 AND Y = 12 else
"000000000000" when X = 73 AND Y = 12 else
"000000000000" when X = 74 AND Y = 12 else
"000000000000" when X = 0 AND Y = 13 else
"000000000000" when X = 1 AND Y = 13 else
"000000000000" when X = 2 AND Y = 13 else
"000000000000" when X = 3 AND Y = 13 else
"000000000000" when X = 4 AND Y = 13 else
"001000100011" when X = 5 AND Y = 13 else
"010101011000" when X = 6 AND Y = 13 else
"100010011101" when X = 7 AND Y = 13 else
"100110101110" when X = 8 AND Y = 13 else
"110011001110" when X = 9 AND Y = 13 else
"110111011111" when X = 10 AND Y = 13 else
"110111011111" when X = 11 AND Y = 13 else
"110111011111" when X = 12 AND Y = 13 else
"110111011111" when X = 13 AND Y = 13 else
"110111011111" when X = 14 AND Y = 13 else
"110111011111" when X = 15 AND Y = 13 else
"110111011111" when X = 16 AND Y = 13 else
"110111011111" when X = 17 AND Y = 13 else
"110111011111" when X = 18 AND Y = 13 else
"110111011111" when X = 19 AND Y = 13 else
"110111011111" when X = 20 AND Y = 13 else
"110111011111" when X = 21 AND Y = 13 else
"111111111111" when X = 22 AND Y = 13 else
"111111111111" when X = 23 AND Y = 13 else
"111111111111" when X = 24 AND Y = 13 else
"111111111111" when X = 25 AND Y = 13 else
"111111111111" when X = 26 AND Y = 13 else
"111111111111" when X = 27 AND Y = 13 else
"111111111111" when X = 28 AND Y = 13 else
"111111111111" when X = 29 AND Y = 13 else
"111111111111" when X = 30 AND Y = 13 else
"111111111111" when X = 31 AND Y = 13 else
"111111111111" when X = 32 AND Y = 13 else
"111111111111" when X = 33 AND Y = 13 else
"111111111111" when X = 34 AND Y = 13 else
"111111111111" when X = 35 AND Y = 13 else
"111111111111" when X = 36 AND Y = 13 else
"111111111111" when X = 37 AND Y = 13 else
"111111111111" when X = 38 AND Y = 13 else
"111111111111" when X = 39 AND Y = 13 else
"111111111111" when X = 40 AND Y = 13 else
"111111111111" when X = 41 AND Y = 13 else
"111111111111" when X = 42 AND Y = 13 else
"111111111111" when X = 43 AND Y = 13 else
"111111111111" when X = 44 AND Y = 13 else
"111111111111" when X = 45 AND Y = 13 else
"111111111111" when X = 46 AND Y = 13 else
"111111111111" when X = 47 AND Y = 13 else
"111111111111" when X = 48 AND Y = 13 else
"111111111111" when X = 49 AND Y = 13 else
"111111111111" when X = 50 AND Y = 13 else
"111111111111" when X = 51 AND Y = 13 else
"111111111111" when X = 52 AND Y = 13 else
"111111111111" when X = 53 AND Y = 13 else
"111111111111" when X = 54 AND Y = 13 else
"111111111111" when X = 55 AND Y = 13 else
"111111111111" when X = 56 AND Y = 13 else
"111111111111" when X = 57 AND Y = 13 else
"111111111111" when X = 58 AND Y = 13 else
"111111111111" when X = 59 AND Y = 13 else
"111111111111" when X = 60 AND Y = 13 else
"110111101111" when X = 61 AND Y = 13 else
"110111011111" when X = 62 AND Y = 13 else
"110111011111" when X = 63 AND Y = 13 else
"101010101100" when X = 64 AND Y = 13 else
"000000000000" when X = 65 AND Y = 13 else
"000000000000" when X = 66 AND Y = 13 else
"000000000000" when X = 67 AND Y = 13 else
"000000000000" when X = 68 AND Y = 13 else
"000000000000" when X = 69 AND Y = 13 else
"000000000000" when X = 70 AND Y = 13 else
"000000000000" when X = 71 AND Y = 13 else
"000000000000" when X = 72 AND Y = 13 else
"000000000000" when X = 73 AND Y = 13 else
"000000000000" when X = 74 AND Y = 13 else
"000000000000" when X = 0 AND Y = 14 else
"000000000000" when X = 1 AND Y = 14 else
"000000000000" when X = 2 AND Y = 14 else
"000000000000" when X = 3 AND Y = 14 else
"001000100011" when X = 4 AND Y = 14 else
"010101011000" when X = 5 AND Y = 14 else
"011110011101" when X = 6 AND Y = 14 else
"100010011101" when X = 7 AND Y = 14 else
"110011001110" when X = 8 AND Y = 14 else
"110111011111" when X = 9 AND Y = 14 else
"110111011111" when X = 10 AND Y = 14 else
"110111011111" when X = 11 AND Y = 14 else
"110111011111" when X = 12 AND Y = 14 else
"110111011111" when X = 13 AND Y = 14 else
"110111011111" when X = 14 AND Y = 14 else
"110111011111" when X = 15 AND Y = 14 else
"110111011111" when X = 16 AND Y = 14 else
"110111011111" when X = 17 AND Y = 14 else
"110111011111" when X = 18 AND Y = 14 else
"110111011111" when X = 19 AND Y = 14 else
"110111011111" when X = 20 AND Y = 14 else
"110111011111" when X = 21 AND Y = 14 else
"110111011111" when X = 22 AND Y = 14 else
"111111111111" when X = 23 AND Y = 14 else
"111111111111" when X = 24 AND Y = 14 else
"111111111111" when X = 25 AND Y = 14 else
"111111111111" when X = 26 AND Y = 14 else
"111111111111" when X = 27 AND Y = 14 else
"111111111111" when X = 28 AND Y = 14 else
"111111111111" when X = 29 AND Y = 14 else
"111111111111" when X = 30 AND Y = 14 else
"111111111111" when X = 31 AND Y = 14 else
"111111111111" when X = 32 AND Y = 14 else
"111111111111" when X = 33 AND Y = 14 else
"111111111111" when X = 34 AND Y = 14 else
"111111111111" when X = 35 AND Y = 14 else
"111111111111" when X = 36 AND Y = 14 else
"111111111111" when X = 37 AND Y = 14 else
"111111111111" when X = 38 AND Y = 14 else
"111111111111" when X = 39 AND Y = 14 else
"111111111111" when X = 40 AND Y = 14 else
"111111111111" when X = 41 AND Y = 14 else
"111111111111" when X = 42 AND Y = 14 else
"111111111111" when X = 43 AND Y = 14 else
"111111111111" when X = 44 AND Y = 14 else
"111111111111" when X = 45 AND Y = 14 else
"111111111111" when X = 46 AND Y = 14 else
"111111111111" when X = 47 AND Y = 14 else
"111111111111" when X = 48 AND Y = 14 else
"111111111111" when X = 49 AND Y = 14 else
"111111111111" when X = 50 AND Y = 14 else
"111111111111" when X = 51 AND Y = 14 else
"111111111111" when X = 52 AND Y = 14 else
"111111111111" when X = 53 AND Y = 14 else
"111111111111" when X = 54 AND Y = 14 else
"111111111111" when X = 55 AND Y = 14 else
"111111111111" when X = 56 AND Y = 14 else
"111111111111" when X = 57 AND Y = 14 else
"111111111111" when X = 58 AND Y = 14 else
"111111111111" when X = 59 AND Y = 14 else
"111111111111" when X = 60 AND Y = 14 else
"110111101111" when X = 61 AND Y = 14 else
"110111011111" when X = 62 AND Y = 14 else
"110111011111" when X = 63 AND Y = 14 else
"101010101100" when X = 64 AND Y = 14 else
"000000000000" when X = 65 AND Y = 14 else
"000000000000" when X = 66 AND Y = 14 else
"000000000000" when X = 67 AND Y = 14 else
"000000000000" when X = 68 AND Y = 14 else
"000000000000" when X = 69 AND Y = 14 else
"000000000000" when X = 70 AND Y = 14 else
"000000000000" when X = 71 AND Y = 14 else
"000000000000" when X = 72 AND Y = 14 else
"000000000000" when X = 73 AND Y = 14 else
"000000000000" when X = 74 AND Y = 14 else
"000000000000" when X = 0 AND Y = 15 else
"000000000000" when X = 1 AND Y = 15 else
"000100100011" when X = 2 AND Y = 15 else
"001000100100" when X = 3 AND Y = 15 else
"010101101001" when X = 4 AND Y = 15 else
"011110001101" when X = 5 AND Y = 15 else
"100010011101" when X = 6 AND Y = 15 else
"100010011101" when X = 7 AND Y = 15 else
"110011011110" when X = 8 AND Y = 15 else
"110111011111" when X = 9 AND Y = 15 else
"110111011111" when X = 10 AND Y = 15 else
"110111011111" when X = 11 AND Y = 15 else
"110111011111" when X = 12 AND Y = 15 else
"110111011111" when X = 13 AND Y = 15 else
"110111011111" when X = 14 AND Y = 15 else
"110111011111" when X = 15 AND Y = 15 else
"110111011111" when X = 16 AND Y = 15 else
"110111011111" when X = 17 AND Y = 15 else
"110111011111" when X = 18 AND Y = 15 else
"110111011111" when X = 19 AND Y = 15 else
"110111011111" when X = 20 AND Y = 15 else
"110111011111" when X = 21 AND Y = 15 else
"110111011111" when X = 22 AND Y = 15 else
"110111011111" when X = 23 AND Y = 15 else
"111111111111" when X = 24 AND Y = 15 else
"111111111111" when X = 25 AND Y = 15 else
"111111111111" when X = 26 AND Y = 15 else
"111111111111" when X = 27 AND Y = 15 else
"111111111111" when X = 28 AND Y = 15 else
"111111111111" when X = 29 AND Y = 15 else
"111111111111" when X = 30 AND Y = 15 else
"111111111111" when X = 31 AND Y = 15 else
"111111111111" when X = 32 AND Y = 15 else
"111111111111" when X = 33 AND Y = 15 else
"111111111111" when X = 34 AND Y = 15 else
"111111111111" when X = 35 AND Y = 15 else
"111111111111" when X = 36 AND Y = 15 else
"111111111111" when X = 37 AND Y = 15 else
"111111111111" when X = 38 AND Y = 15 else
"111111111111" when X = 39 AND Y = 15 else
"111111111111" when X = 40 AND Y = 15 else
"111111111111" when X = 41 AND Y = 15 else
"111111111111" when X = 42 AND Y = 15 else
"111111111111" when X = 43 AND Y = 15 else
"111111111111" when X = 44 AND Y = 15 else
"111111111111" when X = 45 AND Y = 15 else
"111111111111" when X = 46 AND Y = 15 else
"111111111111" when X = 47 AND Y = 15 else
"111111111111" when X = 48 AND Y = 15 else
"111111111111" when X = 49 AND Y = 15 else
"111111111111" when X = 50 AND Y = 15 else
"111111111111" when X = 51 AND Y = 15 else
"111111111111" when X = 52 AND Y = 15 else
"111111111111" when X = 53 AND Y = 15 else
"111111111111" when X = 54 AND Y = 15 else
"111111111111" when X = 55 AND Y = 15 else
"111111111111" when X = 56 AND Y = 15 else
"111111111111" when X = 57 AND Y = 15 else
"111111111111" when X = 58 AND Y = 15 else
"111111111111" when X = 59 AND Y = 15 else
"111111111111" when X = 60 AND Y = 15 else
"110111101111" when X = 61 AND Y = 15 else
"110111011111" when X = 62 AND Y = 15 else
"110111011111" when X = 63 AND Y = 15 else
"101010101100" when X = 64 AND Y = 15 else
"000000000000" when X = 65 AND Y = 15 else
"000000000000" when X = 66 AND Y = 15 else
"000000000000" when X = 67 AND Y = 15 else
"000000000000" when X = 68 AND Y = 15 else
"000000000000" when X = 69 AND Y = 15 else
"000000000000" when X = 70 AND Y = 15 else
"000000000000" when X = 71 AND Y = 15 else
"000000000000" when X = 72 AND Y = 15 else
"000000000000" when X = 73 AND Y = 15 else
"000000000000" when X = 74 AND Y = 15 else
"000000000000" when X = 0 AND Y = 16 else
"000100010010" when X = 1 AND Y = 16 else
"011001111010" when X = 2 AND Y = 16 else
"011110001100" when X = 3 AND Y = 16 else
"011110001101" when X = 4 AND Y = 16 else
"100010011101" when X = 5 AND Y = 16 else
"100010011101" when X = 6 AND Y = 16 else
"110011001110" when X = 7 AND Y = 16 else
"110111011111" when X = 8 AND Y = 16 else
"110111011111" when X = 9 AND Y = 16 else
"110111011111" when X = 10 AND Y = 16 else
"110111011111" when X = 11 AND Y = 16 else
"110111011111" when X = 12 AND Y = 16 else
"110111011111" when X = 13 AND Y = 16 else
"110111011111" when X = 14 AND Y = 16 else
"110111011111" when X = 15 AND Y = 16 else
"110111011111" when X = 16 AND Y = 16 else
"110111011111" when X = 17 AND Y = 16 else
"110111011111" when X = 18 AND Y = 16 else
"110111011111" when X = 19 AND Y = 16 else
"110111011111" when X = 20 AND Y = 16 else
"110111011111" when X = 21 AND Y = 16 else
"110111011111" when X = 22 AND Y = 16 else
"110111011111" when X = 23 AND Y = 16 else
"111111111111" when X = 24 AND Y = 16 else
"111111111111" when X = 25 AND Y = 16 else
"111111111111" when X = 26 AND Y = 16 else
"111111111111" when X = 27 AND Y = 16 else
"111111111111" when X = 28 AND Y = 16 else
"111111111111" when X = 29 AND Y = 16 else
"111111111111" when X = 30 AND Y = 16 else
"111111111111" when X = 31 AND Y = 16 else
"111111111111" when X = 32 AND Y = 16 else
"111111111111" when X = 33 AND Y = 16 else
"111111111111" when X = 34 AND Y = 16 else
"111111111111" when X = 35 AND Y = 16 else
"111111111111" when X = 36 AND Y = 16 else
"111111111111" when X = 37 AND Y = 16 else
"111111111111" when X = 38 AND Y = 16 else
"111111111111" when X = 39 AND Y = 16 else
"111111111111" when X = 40 AND Y = 16 else
"111111111111" when X = 41 AND Y = 16 else
"111111111111" when X = 42 AND Y = 16 else
"111111111111" when X = 43 AND Y = 16 else
"111111111111" when X = 44 AND Y = 16 else
"111111111111" when X = 45 AND Y = 16 else
"111111111111" when X = 46 AND Y = 16 else
"111111111111" when X = 47 AND Y = 16 else
"111111111111" when X = 48 AND Y = 16 else
"111111111111" when X = 49 AND Y = 16 else
"111111111111" when X = 50 AND Y = 16 else
"111111111111" when X = 51 AND Y = 16 else
"111111111111" when X = 52 AND Y = 16 else
"111111111111" when X = 53 AND Y = 16 else
"111111111111" when X = 54 AND Y = 16 else
"111111111111" when X = 55 AND Y = 16 else
"111111111111" when X = 56 AND Y = 16 else
"111111111111" when X = 57 AND Y = 16 else
"111111111111" when X = 58 AND Y = 16 else
"111111111111" when X = 59 AND Y = 16 else
"111111111111" when X = 60 AND Y = 16 else
"110111101111" when X = 61 AND Y = 16 else
"110111011111" when X = 62 AND Y = 16 else
"110111011110" when X = 63 AND Y = 16 else
"101010101011" when X = 64 AND Y = 16 else
"000000000000" when X = 65 AND Y = 16 else
"000000000000" when X = 66 AND Y = 16 else
"000000000000" when X = 67 AND Y = 16 else
"000000000000" when X = 68 AND Y = 16 else
"000000000000" when X = 69 AND Y = 16 else
"000000000000" when X = 70 AND Y = 16 else
"000000000000" when X = 71 AND Y = 16 else
"000000000000" when X = 72 AND Y = 16 else
"000000000000" when X = 73 AND Y = 16 else
"000000000000" when X = 74 AND Y = 16 else
"000100010010" when X = 0 AND Y = 17 else
"011001111010" when X = 1 AND Y = 17 else
"011110001101" when X = 2 AND Y = 17 else
"100010011101" when X = 3 AND Y = 17 else
"100010011101" when X = 4 AND Y = 17 else
"100010011101" when X = 5 AND Y = 17 else
"100110011101" when X = 6 AND Y = 17 else
"110111011110" when X = 7 AND Y = 17 else
"110111011111" when X = 8 AND Y = 17 else
"110111011111" when X = 9 AND Y = 17 else
"110111011111" when X = 10 AND Y = 17 else
"110111011111" when X = 11 AND Y = 17 else
"110111011111" when X = 12 AND Y = 17 else
"110111011111" when X = 13 AND Y = 17 else
"110111011111" when X = 14 AND Y = 17 else
"110111011111" when X = 15 AND Y = 17 else
"110111011111" when X = 16 AND Y = 17 else
"110111011111" when X = 17 AND Y = 17 else
"110111011111" when X = 18 AND Y = 17 else
"110111011111" when X = 19 AND Y = 17 else
"110111011111" when X = 20 AND Y = 17 else
"110111011111" when X = 21 AND Y = 17 else
"110111011111" when X = 22 AND Y = 17 else
"110111011111" when X = 23 AND Y = 17 else
"110111101111" when X = 24 AND Y = 17 else
"111111111111" when X = 25 AND Y = 17 else
"111111111111" when X = 26 AND Y = 17 else
"111111111111" when X = 27 AND Y = 17 else
"111111111111" when X = 28 AND Y = 17 else
"111111111111" when X = 29 AND Y = 17 else
"111111111111" when X = 30 AND Y = 17 else
"111111111111" when X = 31 AND Y = 17 else
"111111111111" when X = 32 AND Y = 17 else
"111111111111" when X = 33 AND Y = 17 else
"111111111111" when X = 34 AND Y = 17 else
"111111111111" when X = 35 AND Y = 17 else
"111111111111" when X = 36 AND Y = 17 else
"111111111111" when X = 37 AND Y = 17 else
"111111111111" when X = 38 AND Y = 17 else
"111111111111" when X = 39 AND Y = 17 else
"111111111111" when X = 40 AND Y = 17 else
"111111111111" when X = 41 AND Y = 17 else
"111111111111" when X = 42 AND Y = 17 else
"111111111111" when X = 43 AND Y = 17 else
"111111111111" when X = 44 AND Y = 17 else
"111111111111" when X = 45 AND Y = 17 else
"111111111111" when X = 46 AND Y = 17 else
"111111111111" when X = 47 AND Y = 17 else
"111111111111" when X = 48 AND Y = 17 else
"111111111111" when X = 49 AND Y = 17 else
"111111111111" when X = 50 AND Y = 17 else
"111111111111" when X = 51 AND Y = 17 else
"111111111111" when X = 52 AND Y = 17 else
"111111111111" when X = 53 AND Y = 17 else
"111111111111" when X = 54 AND Y = 17 else
"111111111111" when X = 55 AND Y = 17 else
"111111111111" when X = 56 AND Y = 17 else
"111111111111" when X = 57 AND Y = 17 else
"111111111111" when X = 58 AND Y = 17 else
"111111111111" when X = 59 AND Y = 17 else
"111111111111" when X = 60 AND Y = 17 else
"110111101111" when X = 61 AND Y = 17 else
"110111011111" when X = 62 AND Y = 17 else
"101010101100" when X = 63 AND Y = 17 else
"010101010110" when X = 64 AND Y = 17 else
"000000000000" when X = 65 AND Y = 17 else
"000000000000" when X = 66 AND Y = 17 else
"000000000000" when X = 67 AND Y = 17 else
"000000000000" when X = 68 AND Y = 17 else
"000000000000" when X = 69 AND Y = 17 else
"000000000000" when X = 70 AND Y = 17 else
"000000000000" when X = 71 AND Y = 17 else
"000000000000" when X = 72 AND Y = 17 else
"000000000000" when X = 73 AND Y = 17 else
"000000000000" when X = 74 AND Y = 17 else
"011001111011" when X = 0 AND Y = 18 else
"011110001101" when X = 1 AND Y = 18 else
"100010011101" when X = 2 AND Y = 18 else
"100010011101" when X = 3 AND Y = 18 else
"100010011101" when X = 4 AND Y = 18 else
"100010011101" when X = 5 AND Y = 18 else
"100010011101" when X = 6 AND Y = 18 else
"110011011110" when X = 7 AND Y = 18 else
"110111011111" when X = 8 AND Y = 18 else
"110111011111" when X = 9 AND Y = 18 else
"110111011111" when X = 10 AND Y = 18 else
"110111011111" when X = 11 AND Y = 18 else
"110111011111" when X = 12 AND Y = 18 else
"110111011111" when X = 13 AND Y = 18 else
"110111011111" when X = 14 AND Y = 18 else
"110111011111" when X = 15 AND Y = 18 else
"110111011111" when X = 16 AND Y = 18 else
"110111011111" when X = 17 AND Y = 18 else
"110111011111" when X = 18 AND Y = 18 else
"110111011111" when X = 19 AND Y = 18 else
"110111011111" when X = 20 AND Y = 18 else
"110111011111" when X = 21 AND Y = 18 else
"110111011111" when X = 22 AND Y = 18 else
"110111011111" when X = 23 AND Y = 18 else
"111011101111" when X = 24 AND Y = 18 else
"111111111111" when X = 25 AND Y = 18 else
"111111111111" when X = 26 AND Y = 18 else
"111111111111" when X = 27 AND Y = 18 else
"111111111111" when X = 28 AND Y = 18 else
"111111111111" when X = 29 AND Y = 18 else
"111111111111" when X = 30 AND Y = 18 else
"111111111111" when X = 31 AND Y = 18 else
"111111111111" when X = 32 AND Y = 18 else
"111111111111" when X = 33 AND Y = 18 else
"111111111111" when X = 34 AND Y = 18 else
"111111111111" when X = 35 AND Y = 18 else
"111111111111" when X = 36 AND Y = 18 else
"111111111111" when X = 37 AND Y = 18 else
"111111111111" when X = 38 AND Y = 18 else
"111111111111" when X = 39 AND Y = 18 else
"111111111111" when X = 40 AND Y = 18 else
"111111111111" when X = 41 AND Y = 18 else
"111111111111" when X = 42 AND Y = 18 else
"111111111111" when X = 43 AND Y = 18 else
"111111111111" when X = 44 AND Y = 18 else
"111111111111" when X = 45 AND Y = 18 else
"111111111111" when X = 46 AND Y = 18 else
"111111111111" when X = 47 AND Y = 18 else
"111111111111" when X = 48 AND Y = 18 else
"111111111111" when X = 49 AND Y = 18 else
"111111111111" when X = 50 AND Y = 18 else
"111111111111" when X = 51 AND Y = 18 else
"111111111111" when X = 52 AND Y = 18 else
"111111111111" when X = 53 AND Y = 18 else
"111111111111" when X = 54 AND Y = 18 else
"111111111111" when X = 55 AND Y = 18 else
"111111111111" when X = 56 AND Y = 18 else
"111111111111" when X = 57 AND Y = 18 else
"111111111111" when X = 58 AND Y = 18 else
"111111111111" when X = 59 AND Y = 18 else
"111111111111" when X = 60 AND Y = 18 else
"111111111111" when X = 61 AND Y = 18 else
"110111101111" when X = 62 AND Y = 18 else
"101111001101" when X = 63 AND Y = 18 else
"101010101100" when X = 64 AND Y = 18 else
"100110011010" when X = 65 AND Y = 18 else
"000000000000" when X = 66 AND Y = 18 else
"000000000000" when X = 67 AND Y = 18 else
"000000000000" when X = 68 AND Y = 18 else
"000000000000" when X = 69 AND Y = 18 else
"000000000000" when X = 70 AND Y = 18 else
"000000000000" when X = 71 AND Y = 18 else
"000000000000" when X = 72 AND Y = 18 else
"000000000000" when X = 73 AND Y = 18 else
"000000000000" when X = 74 AND Y = 18 else
"100010011101" when X = 0 AND Y = 19 else
"100010011101" when X = 1 AND Y = 19 else
"100010011101" when X = 2 AND Y = 19 else
"100010011101" when X = 3 AND Y = 19 else
"100010011101" when X = 4 AND Y = 19 else
"100010011101" when X = 5 AND Y = 19 else
"101110111110" when X = 6 AND Y = 19 else
"110111011111" when X = 7 AND Y = 19 else
"110111011111" when X = 8 AND Y = 19 else
"110111011111" when X = 9 AND Y = 19 else
"110111011111" when X = 10 AND Y = 19 else
"110111011111" when X = 11 AND Y = 19 else
"110111011111" when X = 12 AND Y = 19 else
"110111011111" when X = 13 AND Y = 19 else
"110111011111" when X = 14 AND Y = 19 else
"110111011111" when X = 15 AND Y = 19 else
"110111011111" when X = 16 AND Y = 19 else
"110111011111" when X = 17 AND Y = 19 else
"110111011111" when X = 18 AND Y = 19 else
"110111011111" when X = 19 AND Y = 19 else
"110111011111" when X = 20 AND Y = 19 else
"110111011111" when X = 21 AND Y = 19 else
"110111011111" when X = 22 AND Y = 19 else
"111011101111" when X = 23 AND Y = 19 else
"111111111111" when X = 24 AND Y = 19 else
"111111111111" when X = 25 AND Y = 19 else
"111111111111" when X = 26 AND Y = 19 else
"111111111111" when X = 27 AND Y = 19 else
"111111111111" when X = 28 AND Y = 19 else
"111111111111" when X = 29 AND Y = 19 else
"111111111111" when X = 30 AND Y = 19 else
"111111111111" when X = 31 AND Y = 19 else
"111111111111" when X = 32 AND Y = 19 else
"111111111111" when X = 33 AND Y = 19 else
"111111111111" when X = 34 AND Y = 19 else
"111111111111" when X = 35 AND Y = 19 else
"111111111111" when X = 36 AND Y = 19 else
"111111111111" when X = 37 AND Y = 19 else
"111111111111" when X = 38 AND Y = 19 else
"111111111111" when X = 39 AND Y = 19 else
"111111111111" when X = 40 AND Y = 19 else
"111111111111" when X = 41 AND Y = 19 else
"111111111111" when X = 42 AND Y = 19 else
"111111111111" when X = 43 AND Y = 19 else
"111111111111" when X = 44 AND Y = 19 else
"111111111111" when X = 45 AND Y = 19 else
"111111111111" when X = 46 AND Y = 19 else
"111111111111" when X = 47 AND Y = 19 else
"111111111111" when X = 48 AND Y = 19 else
"111111111111" when X = 49 AND Y = 19 else
"111111111111" when X = 50 AND Y = 19 else
"111111111111" when X = 51 AND Y = 19 else
"111111111111" when X = 52 AND Y = 19 else
"111111111111" when X = 53 AND Y = 19 else
"111111111111" when X = 54 AND Y = 19 else
"111111111111" when X = 55 AND Y = 19 else
"111111111111" when X = 56 AND Y = 19 else
"111111111111" when X = 57 AND Y = 19 else
"111111111111" when X = 58 AND Y = 19 else
"111111111111" when X = 59 AND Y = 19 else
"111111111111" when X = 60 AND Y = 19 else
"111111111111" when X = 61 AND Y = 19 else
"111111111111" when X = 62 AND Y = 19 else
"110111101111" when X = 63 AND Y = 19 else
"110111011111" when X = 64 AND Y = 19 else
"110011001110" when X = 65 AND Y = 19 else
"100110101011" when X = 66 AND Y = 19 else
"100110011010" when X = 67 AND Y = 19 else
"010001000100" when X = 68 AND Y = 19 else
"000000000000" when X = 69 AND Y = 19 else
"000000000000" when X = 70 AND Y = 19 else
"000000000000" when X = 71 AND Y = 19 else
"000000000000" when X = 72 AND Y = 19 else
"000000000000" when X = 73 AND Y = 19 else
"000000000000" when X = 74 AND Y = 19 else
"100010011101" when X = 0 AND Y = 20 else
"100010011101" when X = 1 AND Y = 20 else
"100010011101" when X = 2 AND Y = 20 else
"100010011101" when X = 3 AND Y = 20 else
"100010011101" when X = 4 AND Y = 20 else
"101010111110" when X = 5 AND Y = 20 else
"110111011111" when X = 6 AND Y = 20 else
"110111011111" when X = 7 AND Y = 20 else
"110111011111" when X = 8 AND Y = 20 else
"110111011111" when X = 9 AND Y = 20 else
"110111011111" when X = 10 AND Y = 20 else
"110111011111" when X = 11 AND Y = 20 else
"110111011111" when X = 12 AND Y = 20 else
"110111011111" when X = 13 AND Y = 20 else
"110111011111" when X = 14 AND Y = 20 else
"110111011111" when X = 15 AND Y = 20 else
"111011101111" when X = 16 AND Y = 20 else
"111011101111" when X = 17 AND Y = 20 else
"111011101111" when X = 18 AND Y = 20 else
"111011101111" when X = 19 AND Y = 20 else
"111011101111" when X = 20 AND Y = 20 else
"111011101111" when X = 21 AND Y = 20 else
"111011101111" when X = 22 AND Y = 20 else
"111111111111" when X = 23 AND Y = 20 else
"111111111111" when X = 24 AND Y = 20 else
"111111111111" when X = 25 AND Y = 20 else
"111111111111" when X = 26 AND Y = 20 else
"111111111111" when X = 27 AND Y = 20 else
"111111111111" when X = 28 AND Y = 20 else
"111111111111" when X = 29 AND Y = 20 else
"111111111111" when X = 30 AND Y = 20 else
"111111111111" when X = 31 AND Y = 20 else
"111111111111" when X = 32 AND Y = 20 else
"111111111111" when X = 33 AND Y = 20 else
"111111111111" when X = 34 AND Y = 20 else
"111111111111" when X = 35 AND Y = 20 else
"111111111111" when X = 36 AND Y = 20 else
"111111111111" when X = 37 AND Y = 20 else
"111111111111" when X = 38 AND Y = 20 else
"111111111111" when X = 39 AND Y = 20 else
"111111111111" when X = 40 AND Y = 20 else
"111111111111" when X = 41 AND Y = 20 else
"111111111111" when X = 42 AND Y = 20 else
"111111111111" when X = 43 AND Y = 20 else
"111111111111" when X = 44 AND Y = 20 else
"111111111111" when X = 45 AND Y = 20 else
"111111111111" when X = 46 AND Y = 20 else
"111111111111" when X = 47 AND Y = 20 else
"111111111111" when X = 48 AND Y = 20 else
"111111111111" when X = 49 AND Y = 20 else
"111111111111" when X = 50 AND Y = 20 else
"111111111111" when X = 51 AND Y = 20 else
"111111111111" when X = 52 AND Y = 20 else
"111111111111" when X = 53 AND Y = 20 else
"111111111111" when X = 54 AND Y = 20 else
"111111111111" when X = 55 AND Y = 20 else
"111111111111" when X = 56 AND Y = 20 else
"111111111111" when X = 57 AND Y = 20 else
"111111111111" when X = 58 AND Y = 20 else
"111111111111" when X = 59 AND Y = 20 else
"111111111111" when X = 60 AND Y = 20 else
"111111111111" when X = 61 AND Y = 20 else
"111111111111" when X = 62 AND Y = 20 else
"111011101111" when X = 63 AND Y = 20 else
"110111011111" when X = 64 AND Y = 20 else
"110111011111" when X = 65 AND Y = 20 else
"110111011111" when X = 66 AND Y = 20 else
"110011011110" when X = 67 AND Y = 20 else
"010101010110" when X = 68 AND Y = 20 else
"000000000000" when X = 69 AND Y = 20 else
"000000000000" when X = 70 AND Y = 20 else
"000000000000" when X = 71 AND Y = 20 else
"000000000000" when X = 72 AND Y = 20 else
"000000000000" when X = 73 AND Y = 20 else
"000000000000" when X = 74 AND Y = 20 else
"100010011101" when X = 0 AND Y = 21 else
"100010011101" when X = 1 AND Y = 21 else
"100010011101" when X = 2 AND Y = 21 else
"100010011101" when X = 3 AND Y = 21 else
"101110111110" when X = 4 AND Y = 21 else
"110111011111" when X = 5 AND Y = 21 else
"110111011111" when X = 6 AND Y = 21 else
"110111011111" when X = 7 AND Y = 21 else
"110111011111" when X = 8 AND Y = 21 else
"110111011111" when X = 9 AND Y = 21 else
"110111011111" when X = 10 AND Y = 21 else
"110111011111" when X = 11 AND Y = 21 else
"110111011111" when X = 12 AND Y = 21 else
"110111011111" when X = 13 AND Y = 21 else
"110111011111" when X = 14 AND Y = 21 else
"110111011111" when X = 15 AND Y = 21 else
"111111111111" when X = 16 AND Y = 21 else
"111111111111" when X = 17 AND Y = 21 else
"111111111111" when X = 18 AND Y = 21 else
"111111111111" when X = 19 AND Y = 21 else
"111111111111" when X = 20 AND Y = 21 else
"111111111111" when X = 21 AND Y = 21 else
"111111111111" when X = 22 AND Y = 21 else
"111111111111" when X = 23 AND Y = 21 else
"111111111111" when X = 24 AND Y = 21 else
"111111111111" when X = 25 AND Y = 21 else
"111111111111" when X = 26 AND Y = 21 else
"111111111111" when X = 27 AND Y = 21 else
"111111111111" when X = 28 AND Y = 21 else
"111111111111" when X = 29 AND Y = 21 else
"111111111111" when X = 30 AND Y = 21 else
"111111111111" when X = 31 AND Y = 21 else
"111111111111" when X = 32 AND Y = 21 else
"111111111111" when X = 33 AND Y = 21 else
"111111111111" when X = 34 AND Y = 21 else
"111111111111" when X = 35 AND Y = 21 else
"111111111111" when X = 36 AND Y = 21 else
"111111111111" when X = 37 AND Y = 21 else
"111111111111" when X = 38 AND Y = 21 else
"111111111111" when X = 39 AND Y = 21 else
"111111111111" when X = 40 AND Y = 21 else
"111111111111" when X = 41 AND Y = 21 else
"111111111111" when X = 42 AND Y = 21 else
"111111111111" when X = 43 AND Y = 21 else
"111111111111" when X = 44 AND Y = 21 else
"111111111111" when X = 45 AND Y = 21 else
"111111111111" when X = 46 AND Y = 21 else
"111111111111" when X = 47 AND Y = 21 else
"111111111111" when X = 48 AND Y = 21 else
"111111111111" when X = 49 AND Y = 21 else
"111011111111" when X = 50 AND Y = 21 else
"111011101111" when X = 51 AND Y = 21 else
"111011101111" when X = 52 AND Y = 21 else
"111111111111" when X = 53 AND Y = 21 else
"111111111111" when X = 54 AND Y = 21 else
"111111111111" when X = 55 AND Y = 21 else
"111111111111" when X = 56 AND Y = 21 else
"111111111111" when X = 57 AND Y = 21 else
"111111111111" when X = 58 AND Y = 21 else
"111111111111" when X = 59 AND Y = 21 else
"111111111111" when X = 60 AND Y = 21 else
"111111111111" when X = 61 AND Y = 21 else
"111111111111" when X = 62 AND Y = 21 else
"111011101111" when X = 63 AND Y = 21 else
"110111011111" when X = 64 AND Y = 21 else
"110111011111" when X = 65 AND Y = 21 else
"110111101111" when X = 66 AND Y = 21 else
"110111011110" when X = 67 AND Y = 21 else
"100110011001" when X = 68 AND Y = 21 else
"100010001000" when X = 69 AND Y = 21 else
"011101111000" when X = 70 AND Y = 21 else
"011001110111" when X = 71 AND Y = 21 else
"011001110111" when X = 72 AND Y = 21 else
"011001110111" when X = 73 AND Y = 21 else
"011001110111" when X = 74 AND Y = 21 else
"011110001100" when X = 0 AND Y = 22 else
"100010011101" when X = 1 AND Y = 22 else
"100010011101" when X = 2 AND Y = 22 else
"101010111110" when X = 3 AND Y = 22 else
"110011011110" when X = 4 AND Y = 22 else
"110111011111" when X = 5 AND Y = 22 else
"110111011111" when X = 6 AND Y = 22 else
"110111011111" when X = 7 AND Y = 22 else
"110111011111" when X = 8 AND Y = 22 else
"110111011111" when X = 9 AND Y = 22 else
"110111011111" when X = 10 AND Y = 22 else
"110111011111" when X = 11 AND Y = 22 else
"110111011111" when X = 12 AND Y = 22 else
"110111011111" when X = 13 AND Y = 22 else
"110111011111" when X = 14 AND Y = 22 else
"110111011111" when X = 15 AND Y = 22 else
"111111111111" when X = 16 AND Y = 22 else
"111111111111" when X = 17 AND Y = 22 else
"111111111111" when X = 18 AND Y = 22 else
"111111111111" when X = 19 AND Y = 22 else
"111111111111" when X = 20 AND Y = 22 else
"111111111111" when X = 21 AND Y = 22 else
"111111111111" when X = 22 AND Y = 22 else
"111111111111" when X = 23 AND Y = 22 else
"111111111111" when X = 24 AND Y = 22 else
"111111111111" when X = 25 AND Y = 22 else
"111111111111" when X = 26 AND Y = 22 else
"111111111111" when X = 27 AND Y = 22 else
"111111111111" when X = 28 AND Y = 22 else
"111111111111" when X = 29 AND Y = 22 else
"111111111111" when X = 30 AND Y = 22 else
"111111111111" when X = 31 AND Y = 22 else
"111111111111" when X = 32 AND Y = 22 else
"111111111111" when X = 33 AND Y = 22 else
"111111111111" when X = 34 AND Y = 22 else
"111111111111" when X = 35 AND Y = 22 else
"111111111111" when X = 36 AND Y = 22 else
"111111111111" when X = 37 AND Y = 22 else
"111111111111" when X = 38 AND Y = 22 else
"111111111111" when X = 39 AND Y = 22 else
"111111111111" when X = 40 AND Y = 22 else
"111111111111" when X = 41 AND Y = 22 else
"111111111111" when X = 42 AND Y = 22 else
"111111111111" when X = 43 AND Y = 22 else
"111111111111" when X = 44 AND Y = 22 else
"111111111111" when X = 45 AND Y = 22 else
"111111111111" when X = 46 AND Y = 22 else
"111011101111" when X = 47 AND Y = 22 else
"110111011111" when X = 48 AND Y = 22 else
"110111011111" when X = 49 AND Y = 22 else
"111011101111" when X = 50 AND Y = 22 else
"111111111111" when X = 51 AND Y = 22 else
"111111111111" when X = 52 AND Y = 22 else
"111111111111" when X = 53 AND Y = 22 else
"111111111111" when X = 54 AND Y = 22 else
"111111111111" when X = 55 AND Y = 22 else
"111111111111" when X = 56 AND Y = 22 else
"111111111111" when X = 57 AND Y = 22 else
"111111111111" when X = 58 AND Y = 22 else
"111111111111" when X = 59 AND Y = 22 else
"111111111111" when X = 60 AND Y = 22 else
"111111111111" when X = 61 AND Y = 22 else
"111111111111" when X = 62 AND Y = 22 else
"111011101111" when X = 63 AND Y = 22 else
"110111011111" when X = 64 AND Y = 22 else
"111011101111" when X = 65 AND Y = 22 else
"111111111111" when X = 66 AND Y = 22 else
"111111111111" when X = 67 AND Y = 22 else
"111111111111" when X = 68 AND Y = 22 else
"111111111111" when X = 69 AND Y = 22 else
"111011101111" when X = 70 AND Y = 22 else
"110111011110" when X = 71 AND Y = 22 else
"110111011110" when X = 72 AND Y = 22 else
"110111011110" when X = 73 AND Y = 22 else
"110111011110" when X = 74 AND Y = 22 else
"001100110101" when X = 0 AND Y = 23 else
"011110001100" when X = 1 AND Y = 23 else
"100010011101" when X = 2 AND Y = 23 else
"100010011101" when X = 3 AND Y = 23 else
"101010111110" when X = 4 AND Y = 23 else
"110111011111" when X = 5 AND Y = 23 else
"110111011111" when X = 6 AND Y = 23 else
"110111011111" when X = 7 AND Y = 23 else
"110111011111" when X = 8 AND Y = 23 else
"110111011111" when X = 9 AND Y = 23 else
"110111011111" when X = 10 AND Y = 23 else
"110111011111" when X = 11 AND Y = 23 else
"110111011111" when X = 12 AND Y = 23 else
"110111011111" when X = 13 AND Y = 23 else
"110111011111" when X = 14 AND Y = 23 else
"110111011111" when X = 15 AND Y = 23 else
"111111111111" when X = 16 AND Y = 23 else
"111111111111" when X = 17 AND Y = 23 else
"111111111111" when X = 18 AND Y = 23 else
"111111111111" when X = 19 AND Y = 23 else
"111111111111" when X = 20 AND Y = 23 else
"111111111111" when X = 21 AND Y = 23 else
"111111111111" when X = 22 AND Y = 23 else
"111111111111" when X = 23 AND Y = 23 else
"111111111111" when X = 24 AND Y = 23 else
"111111111111" when X = 25 AND Y = 23 else
"111111111111" when X = 26 AND Y = 23 else
"111111111111" when X = 27 AND Y = 23 else
"111111111111" when X = 28 AND Y = 23 else
"111111111111" when X = 29 AND Y = 23 else
"111111111111" when X = 30 AND Y = 23 else
"111111111111" when X = 31 AND Y = 23 else
"111111111111" when X = 32 AND Y = 23 else
"111111111111" when X = 33 AND Y = 23 else
"111111111111" when X = 34 AND Y = 23 else
"111111111111" when X = 35 AND Y = 23 else
"111111111111" when X = 36 AND Y = 23 else
"110111101111" when X = 37 AND Y = 23 else
"110111011111" when X = 38 AND Y = 23 else
"110111011111" when X = 39 AND Y = 23 else
"110111011111" when X = 40 AND Y = 23 else
"110111011111" when X = 41 AND Y = 23 else
"110111011111" when X = 42 AND Y = 23 else
"110111011111" when X = 43 AND Y = 23 else
"110111011111" when X = 44 AND Y = 23 else
"110111011111" when X = 45 AND Y = 23 else
"110111011111" when X = 46 AND Y = 23 else
"110111011111" when X = 47 AND Y = 23 else
"110111011111" when X = 48 AND Y = 23 else
"111011101111" when X = 49 AND Y = 23 else
"111111111111" when X = 50 AND Y = 23 else
"111111111111" when X = 51 AND Y = 23 else
"111111111111" when X = 52 AND Y = 23 else
"111111111111" when X = 53 AND Y = 23 else
"111111111111" when X = 54 AND Y = 23 else
"111011101111" when X = 55 AND Y = 23 else
"110111011110" when X = 56 AND Y = 23 else
"111011101111" when X = 57 AND Y = 23 else
"111111111111" when X = 58 AND Y = 23 else
"111111111111" when X = 59 AND Y = 23 else
"111111111111" when X = 60 AND Y = 23 else
"111111111111" when X = 61 AND Y = 23 else
"111111111111" when X = 62 AND Y = 23 else
"111011101111" when X = 63 AND Y = 23 else
"111011101111" when X = 64 AND Y = 23 else
"111111111111" when X = 65 AND Y = 23 else
"111111111111" when X = 66 AND Y = 23 else
"111111111111" when X = 67 AND Y = 23 else
"111111111111" when X = 68 AND Y = 23 else
"111111111111" when X = 69 AND Y = 23 else
"111011101111" when X = 70 AND Y = 23 else
"110111011111" when X = 71 AND Y = 23 else
"110111011111" when X = 72 AND Y = 23 else
"110111011111" when X = 73 AND Y = 23 else
"110111011111" when X = 74 AND Y = 23 else
"000100010011" when X = 0 AND Y = 24 else
"011110001100" when X = 1 AND Y = 24 else
"100010011101" when X = 2 AND Y = 24 else
"100010011101" when X = 3 AND Y = 24 else
"100010011101" when X = 4 AND Y = 24 else
"101010111110" when X = 5 AND Y = 24 else
"110111011111" when X = 6 AND Y = 24 else
"110111011111" when X = 7 AND Y = 24 else
"110111011111" when X = 8 AND Y = 24 else
"110111011111" when X = 9 AND Y = 24 else
"110111011111" when X = 10 AND Y = 24 else
"110111011111" when X = 11 AND Y = 24 else
"110111011111" when X = 12 AND Y = 24 else
"110111011111" when X = 13 AND Y = 24 else
"110111011111" when X = 14 AND Y = 24 else
"110111011111" when X = 15 AND Y = 24 else
"111111111111" when X = 16 AND Y = 24 else
"111111111111" when X = 17 AND Y = 24 else
"111111111111" when X = 18 AND Y = 24 else
"111111111111" when X = 19 AND Y = 24 else
"111111111111" when X = 20 AND Y = 24 else
"111111111111" when X = 21 AND Y = 24 else
"111111111111" when X = 22 AND Y = 24 else
"111111111111" when X = 23 AND Y = 24 else
"111111111111" when X = 24 AND Y = 24 else
"111111111111" when X = 25 AND Y = 24 else
"111111111111" when X = 26 AND Y = 24 else
"111111111111" when X = 27 AND Y = 24 else
"111111111111" when X = 28 AND Y = 24 else
"111111111111" when X = 29 AND Y = 24 else
"111111111111" when X = 30 AND Y = 24 else
"111111111111" when X = 31 AND Y = 24 else
"111111111111" when X = 32 AND Y = 24 else
"111111111111" when X = 33 AND Y = 24 else
"111111111111" when X = 34 AND Y = 24 else
"111111111111" when X = 35 AND Y = 24 else
"111111111111" when X = 36 AND Y = 24 else
"110111011111" when X = 37 AND Y = 24 else
"110111011111" when X = 38 AND Y = 24 else
"110111011111" when X = 39 AND Y = 24 else
"110111011111" when X = 40 AND Y = 24 else
"110111011111" when X = 41 AND Y = 24 else
"110111011111" when X = 42 AND Y = 24 else
"110111011111" when X = 43 AND Y = 24 else
"110111011111" when X = 44 AND Y = 24 else
"110111011111" when X = 45 AND Y = 24 else
"110111011111" when X = 46 AND Y = 24 else
"111011101111" when X = 47 AND Y = 24 else
"111111111111" when X = 48 AND Y = 24 else
"111011101111" when X = 49 AND Y = 24 else
"110111101111" when X = 50 AND Y = 24 else
"110111101111" when X = 51 AND Y = 24 else
"110111101111" when X = 52 AND Y = 24 else
"110111101111" when X = 53 AND Y = 24 else
"110111101111" when X = 54 AND Y = 24 else
"110111011111" when X = 55 AND Y = 24 else
"101010101100" when X = 56 AND Y = 24 else
"100110011010" when X = 57 AND Y = 24 else
"110111101111" when X = 58 AND Y = 24 else
"110111101111" when X = 59 AND Y = 24 else
"110111101111" when X = 60 AND Y = 24 else
"110111101111" when X = 61 AND Y = 24 else
"110111101111" when X = 62 AND Y = 24 else
"110111011111" when X = 63 AND Y = 24 else
"111011101111" when X = 64 AND Y = 24 else
"111111111111" when X = 65 AND Y = 24 else
"111111111111" when X = 66 AND Y = 24 else
"111111111111" when X = 67 AND Y = 24 else
"111111111111" when X = 68 AND Y = 24 else
"111111111111" when X = 69 AND Y = 24 else
"111011101111" when X = 70 AND Y = 24 else
"110111011111" when X = 71 AND Y = 24 else
"110111011111" when X = 72 AND Y = 24 else
"110111011111" when X = 73 AND Y = 24 else
"110111011111" when X = 74 AND Y = 24 else
"000000000001" when X = 0 AND Y = 25 else
"010001000111" when X = 1 AND Y = 25 else
"011110001100" when X = 2 AND Y = 25 else
"100010011101" when X = 3 AND Y = 25 else
"100010011101" when X = 4 AND Y = 25 else
"100110101110" when X = 5 AND Y = 25 else
"110111011111" when X = 6 AND Y = 25 else
"110111011111" when X = 7 AND Y = 25 else
"110111011111" when X = 8 AND Y = 25 else
"110111011111" when X = 9 AND Y = 25 else
"110111011111" when X = 10 AND Y = 25 else
"110111011111" when X = 11 AND Y = 25 else
"110111011111" when X = 12 AND Y = 25 else
"110111011111" when X = 13 AND Y = 25 else
"110111011111" when X = 14 AND Y = 25 else
"110111011111" when X = 15 AND Y = 25 else
"111111111111" when X = 16 AND Y = 25 else
"111111111111" when X = 17 AND Y = 25 else
"111111111111" when X = 18 AND Y = 25 else
"111111111111" when X = 19 AND Y = 25 else
"111111111111" when X = 20 AND Y = 25 else
"111111111111" when X = 21 AND Y = 25 else
"111111111111" when X = 22 AND Y = 25 else
"111111111111" when X = 23 AND Y = 25 else
"111111111111" when X = 24 AND Y = 25 else
"111111111111" when X = 25 AND Y = 25 else
"111111111111" when X = 26 AND Y = 25 else
"111111111111" when X = 27 AND Y = 25 else
"111111111111" when X = 28 AND Y = 25 else
"111111111111" when X = 29 AND Y = 25 else
"111111111111" when X = 30 AND Y = 25 else
"111111111111" when X = 31 AND Y = 25 else
"111111111111" when X = 32 AND Y = 25 else
"111111111111" when X = 33 AND Y = 25 else
"111111111111" when X = 34 AND Y = 25 else
"111111111111" when X = 35 AND Y = 25 else
"111111111111" when X = 36 AND Y = 25 else
"111111111111" when X = 37 AND Y = 25 else
"111111111111" when X = 38 AND Y = 25 else
"111111111111" when X = 39 AND Y = 25 else
"111111111111" when X = 40 AND Y = 25 else
"111111111111" when X = 41 AND Y = 25 else
"111111111111" when X = 42 AND Y = 25 else
"111111111111" when X = 43 AND Y = 25 else
"111111111111" when X = 44 AND Y = 25 else
"111111111111" when X = 45 AND Y = 25 else
"111111111111" when X = 46 AND Y = 25 else
"111111111111" when X = 47 AND Y = 25 else
"111111111111" when X = 48 AND Y = 25 else
"110111101111" when X = 49 AND Y = 25 else
"110011001101" when X = 50 AND Y = 25 else
"011110001000" when X = 51 AND Y = 25 else
"011101111000" when X = 52 AND Y = 25 else
"011101111000" when X = 53 AND Y = 25 else
"011101111000" when X = 54 AND Y = 25 else
"011101111000" when X = 55 AND Y = 25 else
"010101010110" when X = 56 AND Y = 25 else
"011110001001" when X = 57 AND Y = 25 else
"110111011111" when X = 58 AND Y = 25 else
"110111011111" when X = 59 AND Y = 25 else
"110111011111" when X = 60 AND Y = 25 else
"110111011111" when X = 61 AND Y = 25 else
"110111011111" when X = 62 AND Y = 25 else
"110111011111" when X = 63 AND Y = 25 else
"111011101111" when X = 64 AND Y = 25 else
"111111111111" when X = 65 AND Y = 25 else
"111111111111" when X = 66 AND Y = 25 else
"111111111111" when X = 67 AND Y = 25 else
"111111111111" when X = 68 AND Y = 25 else
"111111111111" when X = 69 AND Y = 25 else
"111011101111" when X = 70 AND Y = 25 else
"110111011111" when X = 71 AND Y = 25 else
"110111011111" when X = 72 AND Y = 25 else
"110111011111" when X = 73 AND Y = 25 else
"110111011111" when X = 74 AND Y = 25 else
"000000000000" when X = 0 AND Y = 26 else
"000000000000" when X = 1 AND Y = 26 else
"011001111011" when X = 2 AND Y = 26 else
"100010011101" when X = 3 AND Y = 26 else
"100010011101" when X = 4 AND Y = 26 else
"100010011101" when X = 5 AND Y = 26 else
"101010111110" when X = 6 AND Y = 26 else
"110111011111" when X = 7 AND Y = 26 else
"110111011111" when X = 8 AND Y = 26 else
"110111011111" when X = 9 AND Y = 26 else
"110111011111" when X = 10 AND Y = 26 else
"110111011111" when X = 11 AND Y = 26 else
"110111011111" when X = 12 AND Y = 26 else
"110111011111" when X = 13 AND Y = 26 else
"110111011111" when X = 14 AND Y = 26 else
"110111011111" when X = 15 AND Y = 26 else
"111011101111" when X = 16 AND Y = 26 else
"111011101111" when X = 17 AND Y = 26 else
"111011101111" when X = 18 AND Y = 26 else
"111011101111" when X = 19 AND Y = 26 else
"111011101111" when X = 20 AND Y = 26 else
"111011101111" when X = 21 AND Y = 26 else
"111011101111" when X = 22 AND Y = 26 else
"111011101111" when X = 23 AND Y = 26 else
"111011101111" when X = 24 AND Y = 26 else
"111011101111" when X = 25 AND Y = 26 else
"111011101111" when X = 26 AND Y = 26 else
"111011101111" when X = 27 AND Y = 26 else
"111011101111" when X = 28 AND Y = 26 else
"111011101111" when X = 29 AND Y = 26 else
"111011101111" when X = 30 AND Y = 26 else
"111011101111" when X = 31 AND Y = 26 else
"111011101111" when X = 32 AND Y = 26 else
"111111111111" when X = 33 AND Y = 26 else
"111111111111" when X = 34 AND Y = 26 else
"111111111111" when X = 35 AND Y = 26 else
"111111111111" when X = 36 AND Y = 26 else
"111111111111" when X = 37 AND Y = 26 else
"111111111111" when X = 38 AND Y = 26 else
"111111111111" when X = 39 AND Y = 26 else
"111111111111" when X = 40 AND Y = 26 else
"111111111111" when X = 41 AND Y = 26 else
"111111111111" when X = 42 AND Y = 26 else
"111111111111" when X = 43 AND Y = 26 else
"111111111111" when X = 44 AND Y = 26 else
"111111111111" when X = 45 AND Y = 26 else
"111111111111" when X = 46 AND Y = 26 else
"111111111111" when X = 47 AND Y = 26 else
"110111101111" when X = 48 AND Y = 26 else
"110111011111" when X = 49 AND Y = 26 else
"101110111101" when X = 50 AND Y = 26 else
"000100010001" when X = 51 AND Y = 26 else
"000000000000" when X = 52 AND Y = 26 else
"000000000000" when X = 53 AND Y = 26 else
"000000000000" when X = 54 AND Y = 26 else
"000000000000" when X = 55 AND Y = 26 else
"000000000000" when X = 56 AND Y = 26 else
"100010001001" when X = 57 AND Y = 26 else
"110111011111" when X = 58 AND Y = 26 else
"110111011111" when X = 59 AND Y = 26 else
"110111011111" when X = 60 AND Y = 26 else
"110111011111" when X = 61 AND Y = 26 else
"110111011111" when X = 62 AND Y = 26 else
"110111011111" when X = 63 AND Y = 26 else
"111011101111" when X = 64 AND Y = 26 else
"111111111111" when X = 65 AND Y = 26 else
"111111111111" when X = 66 AND Y = 26 else
"111111111111" when X = 67 AND Y = 26 else
"111111111111" when X = 68 AND Y = 26 else
"111011111111" when X = 69 AND Y = 26 else
"110111101111" when X = 70 AND Y = 26 else
"110111011111" when X = 71 AND Y = 26 else
"110111011111" when X = 72 AND Y = 26 else
"110111011111" when X = 73 AND Y = 26 else
"110111011111" when X = 74 AND Y = 26 else
"000000000000" when X = 0 AND Y = 27 else
"000000000000" when X = 1 AND Y = 27 else
"010101011000" when X = 2 AND Y = 27 else
"011001101010" when X = 3 AND Y = 27 else
"011110001011" when X = 4 AND Y = 27 else
"100010011101" when X = 5 AND Y = 27 else
"100010011101" when X = 6 AND Y = 27 else
"101010111110" when X = 7 AND Y = 27 else
"101110111110" when X = 8 AND Y = 27 else
"110011011110" when X = 9 AND Y = 27 else
"110111011111" when X = 10 AND Y = 27 else
"110111011111" when X = 11 AND Y = 27 else
"110111011111" when X = 12 AND Y = 27 else
"110111011111" when X = 13 AND Y = 27 else
"110111011111" when X = 14 AND Y = 27 else
"110111011111" when X = 15 AND Y = 27 else
"110111011111" when X = 16 AND Y = 27 else
"110111011111" when X = 17 AND Y = 27 else
"110111011111" when X = 18 AND Y = 27 else
"110111011111" when X = 19 AND Y = 27 else
"110111011111" when X = 20 AND Y = 27 else
"110111011111" when X = 21 AND Y = 27 else
"110111011111" when X = 22 AND Y = 27 else
"110111011111" when X = 23 AND Y = 27 else
"110111011111" when X = 24 AND Y = 27 else
"110111011111" when X = 25 AND Y = 27 else
"110111011111" when X = 26 AND Y = 27 else
"110111011111" when X = 27 AND Y = 27 else
"110111011111" when X = 28 AND Y = 27 else
"110111011111" when X = 29 AND Y = 27 else
"110111011111" when X = 30 AND Y = 27 else
"110111011111" when X = 31 AND Y = 27 else
"110111011111" when X = 32 AND Y = 27 else
"111011101111" when X = 33 AND Y = 27 else
"111011101111" when X = 34 AND Y = 27 else
"111011101111" when X = 35 AND Y = 27 else
"111011101111" when X = 36 AND Y = 27 else
"111011111111" when X = 37 AND Y = 27 else
"111111111111" when X = 38 AND Y = 27 else
"111111111111" when X = 39 AND Y = 27 else
"111111111111" when X = 40 AND Y = 27 else
"111111111111" when X = 41 AND Y = 27 else
"111111111111" when X = 42 AND Y = 27 else
"111111111111" when X = 43 AND Y = 27 else
"111011111111" when X = 44 AND Y = 27 else
"111011101111" when X = 45 AND Y = 27 else
"111011101111" when X = 46 AND Y = 27 else
"110111101111" when X = 47 AND Y = 27 else
"110111011111" when X = 48 AND Y = 27 else
"110111011111" when X = 49 AND Y = 27 else
"101111001101" when X = 50 AND Y = 27 else
"001000100010" when X = 51 AND Y = 27 else
"000000000000" when X = 52 AND Y = 27 else
"000000000000" when X = 53 AND Y = 27 else
"000000000000" when X = 54 AND Y = 27 else
"000000000000" when X = 55 AND Y = 27 else
"000000000000" when X = 56 AND Y = 27 else
"011001100111" when X = 57 AND Y = 27 else
"101110111100" when X = 58 AND Y = 27 else
"110111011110" when X = 59 AND Y = 27 else
"110111011111" when X = 60 AND Y = 27 else
"110111011111" when X = 61 AND Y = 27 else
"110111011111" when X = 62 AND Y = 27 else
"110111011111" when X = 63 AND Y = 27 else
"110111101111" when X = 64 AND Y = 27 else
"111011101111" when X = 65 AND Y = 27 else
"111011101111" when X = 66 AND Y = 27 else
"111011101111" when X = 67 AND Y = 27 else
"111011101111" when X = 68 AND Y = 27 else
"110111101111" when X = 69 AND Y = 27 else
"110111011111" when X = 70 AND Y = 27 else
"110111011111" when X = 71 AND Y = 27 else
"110111011111" when X = 72 AND Y = 27 else
"110111011111" when X = 73 AND Y = 27 else
"110111011111" when X = 74 AND Y = 27 else
"000000000000" when X = 0 AND Y = 28 else
"000000000000" when X = 1 AND Y = 28 else
"000000000000" when X = 2 AND Y = 28 else
"000000000000" when X = 3 AND Y = 28 else
"010001000111" when X = 4 AND Y = 28 else
"011001111011" when X = 5 AND Y = 28 else
"011101111011" when X = 6 AND Y = 28 else
"100010011101" when X = 7 AND Y = 28 else
"100010011101" when X = 8 AND Y = 28 else
"101010111110" when X = 9 AND Y = 28 else
"101111001110" when X = 10 AND Y = 28 else
"101111001110" when X = 11 AND Y = 28 else
"101111001110" when X = 12 AND Y = 28 else
"101111001110" when X = 13 AND Y = 28 else
"101111001110" when X = 14 AND Y = 28 else
"101111001110" when X = 15 AND Y = 28 else
"101111001110" when X = 16 AND Y = 28 else
"101111001110" when X = 17 AND Y = 28 else
"101111001110" when X = 18 AND Y = 28 else
"101111001110" when X = 19 AND Y = 28 else
"101111001110" when X = 20 AND Y = 28 else
"101111001110" when X = 21 AND Y = 28 else
"101111001110" when X = 22 AND Y = 28 else
"101110111101" when X = 23 AND Y = 28 else
"101110111100" when X = 24 AND Y = 28 else
"101110111100" when X = 25 AND Y = 28 else
"101110111100" when X = 26 AND Y = 28 else
"101110111100" when X = 27 AND Y = 28 else
"101111001101" when X = 28 AND Y = 28 else
"110111011111" when X = 29 AND Y = 28 else
"110111011111" when X = 30 AND Y = 28 else
"110111011111" when X = 31 AND Y = 28 else
"110111011111" when X = 32 AND Y = 28 else
"110111011111" when X = 33 AND Y = 28 else
"110111011111" when X = 34 AND Y = 28 else
"110111011111" when X = 35 AND Y = 28 else
"110111011111" when X = 36 AND Y = 28 else
"110111011111" when X = 37 AND Y = 28 else
"111011101111" when X = 38 AND Y = 28 else
"111111111111" when X = 39 AND Y = 28 else
"111111111111" when X = 40 AND Y = 28 else
"111111111111" when X = 41 AND Y = 28 else
"111111111111" when X = 42 AND Y = 28 else
"111011101111" when X = 43 AND Y = 28 else
"110111011111" when X = 44 AND Y = 28 else
"110111011111" when X = 45 AND Y = 28 else
"110111011111" when X = 46 AND Y = 28 else
"110111011111" when X = 47 AND Y = 28 else
"110111011111" when X = 48 AND Y = 28 else
"110011001110" when X = 49 AND Y = 28 else
"100110101011" when X = 50 AND Y = 28 else
"000100010001" when X = 51 AND Y = 28 else
"000000000000" when X = 52 AND Y = 28 else
"000000000000" when X = 53 AND Y = 28 else
"000000000000" when X = 54 AND Y = 28 else
"000000000000" when X = 55 AND Y = 28 else
"000000000000" when X = 56 AND Y = 28 else
"000000000000" when X = 57 AND Y = 28 else
"011001100111" when X = 58 AND Y = 28 else
"110111011110" when X = 59 AND Y = 28 else
"110111011111" when X = 60 AND Y = 28 else
"110111011111" when X = 61 AND Y = 28 else
"110111011111" when X = 62 AND Y = 28 else
"110111011111" when X = 63 AND Y = 28 else
"110111011111" when X = 64 AND Y = 28 else
"110011011110" when X = 65 AND Y = 28 else
"101110111100" when X = 66 AND Y = 28 else
"101110111100" when X = 67 AND Y = 28 else
"101110111100" when X = 68 AND Y = 28 else
"101110111100" when X = 69 AND Y = 28 else
"101110111100" when X = 70 AND Y = 28 else
"101110111100" when X = 71 AND Y = 28 else
"101110111100" when X = 72 AND Y = 28 else
"101110111100" when X = 73 AND Y = 28 else
"101110111100" when X = 74 AND Y = 28 else
"000000000000" when X = 0 AND Y = 29 else
"000000000000" when X = 1 AND Y = 29 else
"000000000000" when X = 2 AND Y = 29 else
"000000000000" when X = 3 AND Y = 29 else
"000000000000" when X = 4 AND Y = 29 else
"000000000001" when X = 5 AND Y = 29 else
"001100110101" when X = 6 AND Y = 29 else
"011101111011" when X = 7 AND Y = 29 else
"011110001100" when X = 8 AND Y = 29 else
"100010011101" when X = 9 AND Y = 29 else
"100010011101" when X = 10 AND Y = 29 else
"100010011101" when X = 11 AND Y = 29 else
"100010011101" when X = 12 AND Y = 29 else
"100010011101" when X = 13 AND Y = 29 else
"100010011101" when X = 14 AND Y = 29 else
"100010011101" when X = 15 AND Y = 29 else
"100010011101" when X = 16 AND Y = 29 else
"100010011101" when X = 17 AND Y = 29 else
"100010011101" when X = 18 AND Y = 29 else
"011110001101" when X = 19 AND Y = 29 else
"011110001100" when X = 20 AND Y = 29 else
"011110001100" when X = 21 AND Y = 29 else
"011101111011" when X = 22 AND Y = 29 else
"001100110101" when X = 23 AND Y = 29 else
"000100010001" when X = 24 AND Y = 29 else
"000100010001" when X = 25 AND Y = 29 else
"000100010001" when X = 26 AND Y = 29 else
"000100010001" when X = 27 AND Y = 29 else
"011001100110" when X = 28 AND Y = 29 else
"101111001101" when X = 29 AND Y = 29 else
"110011001101" when X = 30 AND Y = 29 else
"110111011110" when X = 31 AND Y = 29 else
"110111011111" when X = 32 AND Y = 29 else
"110111011111" when X = 33 AND Y = 29 else
"110111011111" when X = 34 AND Y = 29 else
"110111011111" when X = 35 AND Y = 29 else
"110111011111" when X = 36 AND Y = 29 else
"110111011111" when X = 37 AND Y = 29 else
"110111011111" when X = 38 AND Y = 29 else
"110111011111" when X = 39 AND Y = 29 else
"110111011111" when X = 40 AND Y = 29 else
"110111011111" when X = 41 AND Y = 29 else
"110111011111" when X = 42 AND Y = 29 else
"110111011111" when X = 43 AND Y = 29 else
"110111011110" when X = 44 AND Y = 29 else
"110011001101" when X = 45 AND Y = 29 else
"110011001101" when X = 46 AND Y = 29 else
"110011001101" when X = 47 AND Y = 29 else
"110011001101" when X = 48 AND Y = 29 else
"100110011010" when X = 49 AND Y = 29 else
"000100010001" when X = 50 AND Y = 29 else
"000000000000" when X = 51 AND Y = 29 else
"000000000000" when X = 52 AND Y = 29 else
"000000000000" when X = 53 AND Y = 29 else
"000000000000" when X = 54 AND Y = 29 else
"000000000000" when X = 55 AND Y = 29 else
"000000000000" when X = 56 AND Y = 29 else
"000000000000" when X = 57 AND Y = 29 else
"010101100110" when X = 58 AND Y = 29 else
"101111001101" when X = 59 AND Y = 29 else
"110011001101" when X = 60 AND Y = 29 else
"110011001101" when X = 61 AND Y = 29 else
"110011001101" when X = 62 AND Y = 29 else
"110011001101" when X = 63 AND Y = 29 else
"110011001101" when X = 64 AND Y = 29 else
"101010101011" when X = 65 AND Y = 29 else
"001000100010" when X = 66 AND Y = 29 else
"000100010001" when X = 67 AND Y = 29 else
"000100010001" when X = 68 AND Y = 29 else
"000100010001" when X = 69 AND Y = 29 else
"000100010001" when X = 70 AND Y = 29 else
"000100010001" when X = 71 AND Y = 29 else
"000100010001" when X = 72 AND Y = 29 else
"000100010001" when X = 73 AND Y = 29 else
"000100010001" when X = 74 AND Y = 29 else
"000000000000" when X = 0 AND Y = 30 else
"000000000000" when X = 1 AND Y = 30 else
"000000000000" when X = 2 AND Y = 30 else
"000000000000" when X = 3 AND Y = 30 else
"000000000000" when X = 4 AND Y = 30 else
"000000000000" when X = 5 AND Y = 30 else
"000000000001" when X = 6 AND Y = 30 else
"000100100011" when X = 7 AND Y = 30 else
"001000100100" when X = 8 AND Y = 30 else
"011110001011" when X = 9 AND Y = 30 else
"100010011101" when X = 10 AND Y = 30 else
"100010011101" when X = 11 AND Y = 30 else
"100010011101" when X = 12 AND Y = 30 else
"100010011101" when X = 13 AND Y = 30 else
"100010011101" when X = 14 AND Y = 30 else
"100010011101" when X = 15 AND Y = 30 else
"100010011101" when X = 16 AND Y = 30 else
"100010011101" when X = 17 AND Y = 30 else
"100010011101" when X = 18 AND Y = 30 else
"011001111011" when X = 19 AND Y = 30 else
"000100100011" when X = 20 AND Y = 30 else
"000100100011" when X = 21 AND Y = 30 else
"000100100011" when X = 22 AND Y = 30 else
"000000000001" when X = 23 AND Y = 30 else
"000000000000" when X = 24 AND Y = 30 else
"000000000000" when X = 25 AND Y = 30 else
"000000000000" when X = 26 AND Y = 30 else
"000000000000" when X = 27 AND Y = 30 else
"000100010001" when X = 28 AND Y = 30 else
"001100110011" when X = 29 AND Y = 30 else
"010001000101" when X = 30 AND Y = 30 else
"110011001101" when X = 31 AND Y = 30 else
"110111011111" when X = 32 AND Y = 30 else
"110111011111" when X = 33 AND Y = 30 else
"110111011111" when X = 34 AND Y = 30 else
"110111011111" when X = 35 AND Y = 30 else
"110111011111" when X = 36 AND Y = 30 else
"110111011111" when X = 37 AND Y = 30 else
"110111011111" when X = 38 AND Y = 30 else
"110111011111" when X = 39 AND Y = 30 else
"110111011111" when X = 40 AND Y = 30 else
"110111011111" when X = 41 AND Y = 30 else
"110111011111" when X = 42 AND Y = 30 else
"110111011111" when X = 43 AND Y = 30 else
"110011011110" when X = 44 AND Y = 30 else
"010101100110" when X = 45 AND Y = 30 else
"001100110100" when X = 46 AND Y = 30 else
"001100110100" when X = 47 AND Y = 30 else
"001100110100" when X = 48 AND Y = 30 else
"001000100011" when X = 49 AND Y = 30 else
"000000000000" when X = 50 AND Y = 30 else
"000000000000" when X = 51 AND Y = 30 else
"000000000000" when X = 52 AND Y = 30 else
"000000000000" when X = 53 AND Y = 30 else
"000000000000" when X = 54 AND Y = 30 else
"000000000000" when X = 55 AND Y = 30 else
"000000000000" when X = 56 AND Y = 30 else
"000000000000" when X = 57 AND Y = 30 else
"000100010001" when X = 58 AND Y = 30 else
"001100110011" when X = 59 AND Y = 30 else
"001100110100" when X = 60 AND Y = 30 else
"001100110100" when X = 61 AND Y = 30 else
"001100110100" when X = 62 AND Y = 30 else
"001100110100" when X = 63 AND Y = 30 else
"001100110100" when X = 64 AND Y = 30 else
"001100110011" when X = 65 AND Y = 30 else
"000000000000" when X = 66 AND Y = 30 else
"000000000000" when X = 67 AND Y = 30 else
"000000000000" when X = 68 AND Y = 30 else
"000000000000" when X = 69 AND Y = 30 else
"000000000000" when X = 70 AND Y = 30 else
"000000000000" when X = 71 AND Y = 30 else
"000000000000" when X = 72 AND Y = 30 else
"000000000000" when X = 73 AND Y = 30 else
"000000000000" when X = 74 AND Y = 30 else
"000000000000"; -- should never get here
end rtl;
