library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

PACKAGE MY IS
PROCEDURE SQ(SIGNAL Xcur,Ycur,Xpos,Ypos:IN INTEGER;SIGNAL RGB:OUT STD_LOGIC_VECTOR(3 downto 0);SIGNAL DRAW: OUT STD_LOGIC);
PROCEDURE DASH(SIGNAL Xcur,Ycur,Xpos,Ypos:IN INTEGER;SIGNAL RGB:OUT STD_LOGIC_VECTOR(3 downto 0);SIGNAL DRAW: OUT STD_LOGIC);
PROCEDURE SKY(SIGNAL Xcur,Ycur,Xpos,Ypos:IN INTEGER;SIGNAL RGB:OUT STD_LOGIC_VECTOR(3 downto 0);SIGNAL DRAW: OUT STD_LOGIC);
PROCEDURE SKY2(SIGNAL Xcur,Ycur,Xpos,Ypos:IN INTEGER;SIGNAL RGB:OUT STD_LOGIC_VECTOR(3 downto 0);SIGNAL DRAW: OUT STD_LOGIC);
PROCEDURE SKY3(SIGNAL Xcur,Ycur,Xpos,Ypos:IN INTEGER;SIGNAL RGB:OUT STD_LOGIC_VECTOR(3 downto 0);SIGNAL DRAW: OUT STD_LOGIC);
PROCEDURE SKY4(SIGNAL Xcur,Ycur,Xpos,Ypos:IN INTEGER;SIGNAL RGB:OUT STD_LOGIC_VECTOR(3 downto 0);SIGNAL DRAW: OUT STD_LOGIC);
PROCEDURE LINEAR(SIGNAL Xcur,Ycur,X1,Y1,X2,Y2:IN INTEGER;SIGNAL RGB:OUT STD_LOGIC_VECTOR(3 downto 0);SIGNAL DRAW: OUT STD_LOGIC);
PROCEDURE LINEARPOS(SIGNAL Xcur,Ycur,X1,Y1,X2,Y2:IN INTEGER;SIGNAL RGB:OUT STD_LOGIC_VECTOR(3 downto 0);SIGNAL DRAW: OUT STD_LOGIC);
PROCEDURE ROAD(SIGNAL Xcur,Ycur,L1_X1,L1_Y1,L1_X2,L1_Y2,L2_X1,L2_Y1,L2_X2,L2_Y2:IN INTEGER;SIGNAL RGB:OUT STD_LOGIC_VECTOR(3 downto 0);SIGNAL DRAW: OUT STD_LOGIC);
PROCEDURE CAR(SIGNAL Xcur,Ycur,Xpos,Ypos:IN INTEGER;SIGNAL CAR_DATA:IN STD_LOGIC_VECTOR(12 downto 0);SIGNAL RGB:OUT STD_LOGIC_VECTOR(3 downto 0);SIGNAL DRAW: OUT STD_LOGIC);
PROCEDURE CLOUD_PROC(SIGNAL Xcur,Ycur,Xpos,Ypos:IN INTEGER;SIGNAL CLOUD_DATA:IN STD_LOGIC_VECTOR(12 downto 0);SIGNAL RGB:OUT STD_LOGIC_VECTOR(3 downto 0);SIGNAL DRAW: OUT STD_LOGIC);
END MY;

PACKAGE BODY MY IS
PROCEDURE SQ(SIGNAL Xcur,Ycur,Xpos,Ypos:IN INTEGER;SIGNAL RGB:OUT STD_LOGIC_VECTOR(3 downto 0);SIGNAL DRAW: OUT STD_LOGIC) IS
BEGIN
 IF(Xcur>Xpos AND Xcur<(Xpos+1600) AND Ycur>Ypos AND Ycur<(Ypos+1000))THEN
	 RGB<="1111";
	 DRAW<='1';
	 ELSE
	 DRAW<='0';
 END IF;
END SQ;

PROCEDURE DASH(SIGNAL Xcur,Ycur,Xpos,Ypos:IN INTEGER;SIGNAL RGB:OUT STD_LOGIC_VECTOR(3 downto 0);SIGNAL DRAW: OUT STD_LOGIC) IS
BEGIN
 IF(Xcur>Xpos AND Xcur<(Xpos+20) AND Ycur>(Ypos-(Ypos/20)+24) AND Ycur<(Ypos+(Ypos/20)-24)) THEN
	 RGB<="1111";
	 DRAW<='1';
	 ELSE
	 DRAW<='0';
 END IF;
END DASH;

PROCEDURE SKY(SIGNAL Xcur,Ycur,Xpos,Ypos:IN INTEGER;SIGNAL RGB:OUT STD_LOGIC_VECTOR(3 downto 0);SIGNAL DRAW: OUT STD_LOGIC) IS
BEGIN
 IF(Xcur>Xpos AND Xcur<(Xpos+1600) AND Ycur>Ypos AND Ycur<(Ypos+500))THEN
	 RGB<="1111";
	 DRAW<='1';
	 ELSE
	 DRAW<='0';
 END IF;
END SKY;

PROCEDURE SKY2(SIGNAL Xcur,Ycur,Xpos,Ypos:IN INTEGER;SIGNAL RGB:OUT STD_LOGIC_VECTOR(3 downto 0);SIGNAL DRAW: OUT STD_LOGIC) IS
BEGIN
 IF(Xcur>Xpos AND Xcur<(Xpos+1600) AND Ycur>Ypos AND Ycur<(Ypos+425))THEN
	 RGB<="1111";
	 DRAW<='1';
	 ELSE
	 DRAW<='0';
 END IF;
END SKY2;

PROCEDURE SKY3(SIGNAL Xcur,Ycur,Xpos,Ypos:IN INTEGER;SIGNAL RGB:OUT STD_LOGIC_VECTOR(3 downto 0);SIGNAL DRAW: OUT STD_LOGIC) IS
BEGIN
 IF(Xcur>Xpos AND Xcur<(Xpos+1600) AND Ycur>Ypos AND Ycur<(Ypos+375))THEN
	 RGB<="1111";
	 DRAW<='1';
	 ELSE
	 DRAW<='0';
 END IF;
END SKY3;

PROCEDURE SKY4(SIGNAL Xcur,Ycur,Xpos,Ypos:IN INTEGER;SIGNAL RGB:OUT STD_LOGIC_VECTOR(3 downto 0);SIGNAL DRAW: OUT STD_LOGIC) IS
BEGIN
 IF(Xcur>Xpos AND Xcur<(Xpos+1600) AND Ycur>Ypos AND Ycur<(Ypos+350))THEN
	 RGB<="1111";
	 DRAW<='1';
	 ELSE
	 DRAW<='0';
 END IF;
END SKY4;

PROCEDURE LINEAR(SIGNAL Xcur,Ycur,X1,Y1,X2,Y2:IN INTEGER;SIGNAL RGB:OUT STD_LOGIC_VECTOR(3 downto 0);SIGNAL DRAW: OUT STD_LOGIC) IS
BEGIN
 IF (Xcur = ((X2-X1)/(Y2-Y1))*(Ycur - Y1) + X1) AND (Ycur = ((Y2-Y1)/(X2-X1)*(Xcur - X1) + Y1) AND Ycur > Y1 AND Xcur > X1)  THEN
	 RGB<="1111";
	 DRAW<='1';
	 ELSE
	 DRAW<='0';
 END IF;
END LINEAR;

PROCEDURE LINEARPOS(SIGNAL Xcur,Ycur,X1,Y1,X2,Y2:IN INTEGER;SIGNAL RGB:OUT STD_LOGIC_VECTOR(3 downto 0);SIGNAL DRAW: OUT STD_LOGIC) IS
BEGIN
 IF (Xcur = ((X2-X1)/(Y2-Y1))*(Ycur - Y1) + X1) AND (Ycur = ((Y2-Y1)/(X2-X1)*(Xcur - X1) + Y1) AND Ycur > Y1 AND Xcur < X1)  THEN
	 RGB<="1111";
	 DRAW<='1';
	 ELSE
	 DRAW<='0';
 END IF;
END LINEARPOS;

PROCEDURE ROAD(SIGNAL Xcur,Ycur,L1_X1,L1_Y1,L1_X2,L1_Y2,L2_X1,L2_Y1,L2_X2,L2_Y2:IN INTEGER;SIGNAL RGB:OUT STD_LOGIC_VECTOR(3 downto 0);SIGNAL DRAW: OUT STD_LOGIC) IS 
BEGIN
 IF (Xcur > ((L2_X2-L2_X1)/(L2_Y2-L2_Y1))*(Ycur - L2_Y1) + L2_X1) AND (Xcur < ((L1_X2-L1_X1)/(L1_Y2-L1_Y1))*(Ycur - L1_Y1) + L1_X1) AND (Ycur > 500) THEN
	 RGB<="1111";
	 DRAW<='1';
	 ELSE
	 DRAW<='0';
 END IF;
END ROAD;

PROCEDURE CAR(SIGNAL Xcur,Ycur,Xpos,Ypos:IN INTEGER;SIGNAL CAR_DATA:IN STD_LOGIC_VECTOR(12 downto 0);SIGNAL RGB:OUT STD_LOGIC_VECTOR(3 downto 0);SIGNAL DRAW: OUT STD_LOGIC) IS
BEGIN
 IF(Xcur>Xpos AND Xcur<(Xpos+46) AND Ycur>Ypos AND Ycur<(Ypos+30) AND CAR_DATA(0) = '1')  THEN
	 RGB<="1111";
	 DRAW<='1';
	 ELSE
	 DRAW<='0';
 END IF;
END CAR;

PROCEDURE CLOUD_PROC(SIGNAL Xcur,Ycur,Xpos,Ypos:IN INTEGER;SIGNAL CLOUD_DATA:IN STD_LOGIC_VECTOR(12 downto 0);SIGNAL RGB:OUT STD_LOGIC_VECTOR(3 downto 0);SIGNAL DRAW: OUT STD_LOGIC) IS
BEGIN
 IF(Xcur>Xpos AND Xcur<(Xpos+75) AND Ycur>Ypos AND Ycur<(Ypos+31) AND CLOUD_DATA(0) = '1')  THEN
	 RGB<="1111";
	 DRAW<='1';
	 ELSE
	 DRAW<='0';
 END IF;
END CLOUD_PROC;

END MY;